`define IN_DATA(index) in_data``index
`define TEMP_ODD(index) temp_odd``index
`define TEMP_EVEN(index) temp_even``index

module Bubble_Sort(
	clk,
	rst_n,
	in_valid,
	in_data,
	out_valid,
	out_data
	);

input             clk;
input             rst_n;
input             in_valid;
input       [7:0] in_data;
output reg	      out_valid;
output reg	[7:0] out_data;

/*
 * Memory to store in data
*/
reg			[7:0] in_data1;
reg			[7:0] in_data2;
reg			[7:0] in_data3;
reg			[7:0] in_data4;
reg			[7:0] in_data5;
reg			[7:0] in_data6;
reg			[7:0] in_data7;
reg			[7:0] in_data8;
reg			[7:0] in_data9;
reg			[7:0] in_data10;
reg			[7:0] in_data11;
reg			[7:0] in_data12;
reg			[7:0] in_data13;
reg			[7:0] in_data14;
reg			[7:0] in_data15;
reg			[7:0] in_data16;
reg			[7:0] in_data17;
reg			[7:0] in_data18;
reg			[7:0] in_data19;
reg			[7:0] in_data20;
reg			[7:0] in_data21;
reg			[7:0] in_data22;
reg			[7:0] in_data23;
reg			[7:0] in_data24;
reg			[7:0] in_data25;
reg			[7:0] in_data26;
reg			[7:0] in_data27;
reg			[7:0] in_data28;
reg			[7:0] in_data29;
reg			[7:0] in_data30;
reg			[7:0] in_data31;
reg			[7:0] in_data32;
reg			[7:0] in_data33;
reg			[7:0] in_data34;
reg			[7:0] in_data35;
reg			[7:0] in_data36;
reg			[7:0] in_data37;
reg			[7:0] in_data38;
reg			[7:0] in_data39;
reg			[7:0] in_data40;
reg			[7:0] in_data41;
reg			[7:0] in_data42;
reg			[7:0] in_data43;
reg			[7:0] in_data44;
reg			[7:0] in_data45;
reg			[7:0] in_data46;
reg			[7:0] in_data47;
reg			[7:0] in_data48;
reg			[7:0] in_data49;
reg			[7:0] in_data50;
reg			[7:0] in_data51;
reg			[7:0] in_data52;
reg			[7:0] in_data53;
reg			[7:0] in_data54;
reg			[7:0] in_data55;
reg			[7:0] in_data56;
reg			[7:0] in_data57;
reg			[7:0] in_data58;
reg			[7:0] in_data59;
reg			[7:0] in_data60;
reg			[7:0] in_data61;
reg			[7:0] in_data62;
reg			[7:0] in_data63;
reg			[7:0] in_data64;
reg			[7:0] in_data65;
reg			[7:0] in_data66;
reg			[7:0] in_data67;
reg			[7:0] in_data68;
reg			[7:0] in_data69;
reg			[7:0] in_data70;
reg			[7:0] in_data71;
reg			[7:0] in_data72;
reg			[7:0] in_data73;
reg			[7:0] in_data74;
reg			[7:0] in_data75;
reg			[7:0] in_data76;
reg			[7:0] in_data77;
reg			[7:0] in_data78;
reg			[7:0] in_data79;
reg			[7:0] in_data80;
reg			[7:0] in_data81;
reg			[7:0] in_data82;
reg			[7:0] in_data83;
reg			[7:0] in_data84;
reg			[7:0] in_data85;
reg			[7:0] in_data86;
reg			[7:0] in_data87;
reg			[7:0] in_data88;
reg			[7:0] in_data89;
reg			[7:0] in_data90;
reg			[7:0] in_data91;
reg			[7:0] in_data92;
reg			[7:0] in_data93;
reg			[7:0] in_data94;
reg			[7:0] in_data95;
reg			[7:0] in_data96;
reg			[7:0] in_data97;
reg			[7:0] in_data98;
reg			[7:0] in_data99;
reg			[7:0] in_data100;
reg			[7:0] in_data101;
reg			[7:0] in_data102;
reg			[7:0] in_data103;
reg			[7:0] in_data104;
reg			[7:0] in_data105;
reg			[7:0] in_data106;
reg			[7:0] in_data107;
reg			[7:0] in_data108;
reg			[7:0] in_data109;
reg			[7:0] in_data110;
reg			[7:0] in_data111;
reg			[7:0] in_data112;
reg			[7:0] in_data113;
reg			[7:0] in_data114;
reg			[7:0] in_data115;
reg			[7:0] in_data116;
reg			[7:0] in_data117;
reg			[7:0] in_data118;
reg			[7:0] in_data119;
reg			[7:0] in_data120;
reg			[7:0] in_data121;
reg			[7:0] in_data122;
reg			[7:0] in_data123;
reg			[7:0] in_data124;
reg			[7:0] in_data125;
reg			[7:0] in_data126;
reg			[7:0] in_data127;
reg			[7:0] in_data128;
reg			[7:0] in_data129;
reg			[7:0] in_data130;
reg			[7:0] in_data131;
reg			[7:0] in_data132;
reg			[7:0] in_data133;
reg			[7:0] in_data134;
reg			[7:0] in_data135;
reg			[7:0] in_data136;
reg			[7:0] in_data137;
reg			[7:0] in_data138;
reg			[7:0] in_data139;
reg			[7:0] in_data140;
reg			[7:0] in_data141;
reg			[7:0] in_data142;
reg			[7:0] in_data143;
reg			[7:0] in_data144;
reg			[7:0] in_data145;
reg			[7:0] in_data146;
reg			[7:0] in_data147;
reg			[7:0] in_data148;
reg			[7:0] in_data149;
reg			[7:0] in_data150;
reg			[7:0] in_data151;
reg			[7:0] in_data152;
reg			[7:0] in_data153;
reg			[7:0] in_data154;
reg			[7:0] in_data155;
reg			[7:0] in_data156;
reg			[7:0] in_data157;
reg			[7:0] in_data158;
reg			[7:0] in_data159;
reg			[7:0] in_data160;
reg			[7:0] in_data161;
reg			[7:0] in_data162;
reg			[7:0] in_data163;
reg			[7:0] in_data164;
reg			[7:0] in_data165;
reg			[7:0] in_data166;
reg			[7:0] in_data167;
reg			[7:0] in_data168;
reg			[7:0] in_data169;
reg			[7:0] in_data170;
reg			[7:0] in_data171;
reg			[7:0] in_data172;
reg			[7:0] in_data173;
reg			[7:0] in_data174;
reg			[7:0] in_data175;
reg			[7:0] in_data176;
reg			[7:0] in_data177;
reg			[7:0] in_data178;
reg			[7:0] in_data179;
reg			[7:0] in_data180;
reg			[7:0] in_data181;
reg			[7:0] in_data182;
reg			[7:0] in_data183;
reg			[7:0] in_data184;
reg			[7:0] in_data185;
reg			[7:0] in_data186;
reg			[7:0] in_data187;
reg			[7:0] in_data188;
reg			[7:0] in_data189;
reg			[7:0] in_data190;
reg			[7:0] in_data191;
reg			[7:0] in_data192;
reg			[7:0] in_data193;
reg			[7:0] in_data194;
reg			[7:0] in_data195;
reg			[7:0] in_data196;
reg			[7:0] in_data197;
reg			[7:0] in_data198;
reg			[7:0] in_data199;
reg			[7:0] in_data200;
reg			[7:0] in_data201;
reg			[7:0] in_data202;
reg			[7:0] in_data203;
reg			[7:0] in_data204;
reg			[7:0] in_data205;
reg			[7:0] in_data206;
reg			[7:0] in_data207;
reg			[7:0] in_data208;
reg			[7:0] in_data209;
reg			[7:0] in_data210;
reg			[7:0] in_data211;
reg			[7:0] in_data212;
reg			[7:0] in_data213;
reg			[7:0] in_data214;
reg			[7:0] in_data215;
reg			[7:0] in_data216;
reg			[7:0] in_data217;
reg			[7:0] in_data218;
reg			[7:0] in_data219;
reg			[7:0] in_data220;
reg			[7:0] in_data221;
reg			[7:0] in_data222;
reg			[7:0] in_data223;
reg			[7:0] in_data224;
reg			[7:0] in_data225;
reg			[7:0] in_data226;
reg			[7:0] in_data227;
reg			[7:0] in_data228;
reg			[7:0] in_data229;
reg			[7:0] in_data230;
reg			[7:0] in_data231;
reg			[7:0] in_data232;
reg			[7:0] in_data233;
reg			[7:0] in_data234;
reg			[7:0] in_data235;
reg			[7:0] in_data236;
reg			[7:0] in_data237;
reg			[7:0] in_data238;
reg			[7:0] in_data239;
reg			[7:0] in_data240;
reg			[7:0] in_data241;
reg			[7:0] in_data242;
reg			[7:0] in_data243;
reg			[7:0] in_data244;
reg			[7:0] in_data245;
reg			[7:0] in_data246;
reg			[7:0] in_data247;
reg			[7:0] in_data248;
reg			[7:0] in_data249;
reg			[7:0] in_data250;
reg			[7:0] in_data251;
reg			[7:0] in_data252;
reg			[7:0] in_data253;
reg			[7:0] in_data254;
reg			[7:0] in_data255;

/*
 * Store input into memory
*/
reg			[7:0] input_index;
reg				  in_valid_flag; //so that calculation of bubble sort can start right after in_valid is low
reg				  bubble_start_flag; //indicates the start of bubble sort (combinational)
always @(posedge clk) begin
	if (!rst_n) begin
		input_index <= 'd0;
		in_valid_flag <= 1'b0;
		bubble_start_flag <= 1'b0;
		in_data1 <= 'd0;
		in_data2 <= 'd0;
		in_data3 <= 'd0;
		in_data4 <= 'd0;
		in_data5 <= 'd0;
		in_data6 <= 'd0;
		in_data7 <= 'd0;
		in_data8 <= 'd0;
		in_data9 <= 'd0;
		in_data10 <= 'd0;
		in_data11 <= 'd0;
		in_data12 <= 'd0;
		in_data13 <= 'd0;
		in_data14 <= 'd0;
		in_data15 <= 'd0;
		in_data16 <= 'd0;
		in_data17 <= 'd0;
		in_data18 <= 'd0;
		in_data19 <= 'd0;
		in_data20 <= 'd0;
		in_data21 <= 'd0;
		in_data22 <= 'd0;
		in_data23 <= 'd0;
		in_data24 <= 'd0;
		in_data25 <= 'd0;
		in_data26 <= 'd0;
		in_data27 <= 'd0;
		in_data28 <= 'd0;
		in_data29 <= 'd0;
		in_data30 <= 'd0;
		in_data31 <= 'd0;
		in_data32 <= 'd0;
		in_data33 <= 'd0;
		in_data34 <= 'd0;
		in_data35 <= 'd0;
		in_data36 <= 'd0;
		in_data37 <= 'd0;
		in_data38 <= 'd0;
		in_data39 <= 'd0;
		in_data40 <= 'd0;
		in_data41 <= 'd0;
		in_data42 <= 'd0;
		in_data43 <= 'd0;
		in_data44 <= 'd0;
		in_data45 <= 'd0;
		in_data46 <= 'd0;
		in_data47 <= 'd0;
		in_data48 <= 'd0;
		in_data49 <= 'd0;
		in_data50 <= 'd0;
		in_data51 <= 'd0;
		in_data52 <= 'd0;
		in_data53 <= 'd0;
		in_data54 <= 'd0;
		in_data55 <= 'd0;
		in_data56 <= 'd0;
		in_data57 <= 'd0;
		in_data58 <= 'd0;
		in_data59 <= 'd0;
		in_data60 <= 'd0;
		in_data61 <= 'd0;
		in_data62 <= 'd0;
		in_data63 <= 'd0;
		in_data64 <= 'd0;
		in_data65 <= 'd0;
		in_data66 <= 'd0;
		in_data67 <= 'd0;
		in_data68 <= 'd0;
		in_data69 <= 'd0;
		in_data70 <= 'd0;
		in_data71 <= 'd0;
		in_data72 <= 'd0;
		in_data73 <= 'd0;
		in_data74 <= 'd0;
		in_data75 <= 'd0;
		in_data76 <= 'd0;
		in_data77 <= 'd0;
		in_data78 <= 'd0;
		in_data79 <= 'd0;
		in_data80 <= 'd0;
		in_data81 <= 'd0;
		in_data82 <= 'd0;
		in_data83 <= 'd0;
		in_data84 <= 'd0;
		in_data85 <= 'd0;
		in_data86 <= 'd0;
		in_data87 <= 'd0;
		in_data88 <= 'd0;
		in_data89 <= 'd0;
		in_data90 <= 'd0;
		in_data91 <= 'd0;
		in_data92 <= 'd0;
		in_data93 <= 'd0;
		in_data94 <= 'd0;
		in_data95 <= 'd0;
		in_data96 <= 'd0;
		in_data97 <= 'd0;
		in_data98 <= 'd0;
		in_data99 <= 'd0;
		in_data100 <= 'd0;
		in_data101 <= 'd0;
		in_data102 <= 'd0;
		in_data103 <= 'd0;
		in_data104 <= 'd0;
		in_data105 <= 'd0;
		in_data106 <= 'd0;
		in_data107 <= 'd0;
		in_data108 <= 'd0;
		in_data109 <= 'd0;
		in_data110 <= 'd0;
		in_data111 <= 'd0;
		in_data112 <= 'd0;
		in_data113 <= 'd0;
		in_data114 <= 'd0;
		in_data115 <= 'd0;
		in_data116 <= 'd0;
		in_data117 <= 'd0;
		in_data118 <= 'd0;
		in_data119 <= 'd0;
		in_data120 <= 'd0;
		in_data121 <= 'd0;
		in_data122 <= 'd0;
		in_data123 <= 'd0;
		in_data124 <= 'd0;
		in_data125 <= 'd0;
		in_data126 <= 'd0;
		in_data127 <= 'd0;
		in_data128 <= 'd0;
		in_data129 <= 'd0;
		in_data130 <= 'd0;
		in_data131 <= 'd0;
		in_data132 <= 'd0;
		in_data133 <= 'd0;
		in_data134 <= 'd0;
		in_data135 <= 'd0;
		in_data136 <= 'd0;
		in_data137 <= 'd0;
		in_data138 <= 'd0;
		in_data139 <= 'd0;
		in_data140 <= 'd0;
		in_data141 <= 'd0;
		in_data142 <= 'd0;
		in_data143 <= 'd0;
		in_data144 <= 'd0;
		in_data145 <= 'd0;
		in_data146 <= 'd0;
		in_data147 <= 'd0;
		in_data148 <= 'd0;
		in_data149 <= 'd0;
		in_data150 <= 'd0;
		in_data151 <= 'd0;
		in_data152 <= 'd0;
		in_data153 <= 'd0;
		in_data154 <= 'd0;
		in_data155 <= 'd0;
		in_data156 <= 'd0;
		in_data157 <= 'd0;
		in_data158 <= 'd0;
		in_data159 <= 'd0;
		in_data160 <= 'd0;
		in_data161 <= 'd0;
		in_data162 <= 'd0;
		in_data163 <= 'd0;
		in_data164 <= 'd0;
		in_data165 <= 'd0;
		in_data166 <= 'd0;
		in_data167 <= 'd0;
		in_data168 <= 'd0;
		in_data169 <= 'd0;
		in_data170 <= 'd0;
		in_data171 <= 'd0;
		in_data172 <= 'd0;
		in_data173 <= 'd0;
		in_data174 <= 'd0;
		in_data175 <= 'd0;
		in_data176 <= 'd0;
		in_data177 <= 'd0;
		in_data178 <= 'd0;
		in_data179 <= 'd0;
		in_data180 <= 'd0;
		in_data181 <= 'd0;
		in_data182 <= 'd0;
		in_data183 <= 'd0;
		in_data184 <= 'd0;
		in_data185 <= 'd0;
		in_data186 <= 'd0;
		in_data187 <= 'd0;
		in_data188 <= 'd0;
		in_data189 <= 'd0;
		in_data190 <= 'd0;
		in_data191 <= 'd0;
		in_data192 <= 'd0;
		in_data193 <= 'd0;
		in_data194 <= 'd0;
		in_data195 <= 'd0;
		in_data196 <= 'd0;
		in_data197 <= 'd0;
		in_data198 <= 'd0;
		in_data199 <= 'd0;
		in_data200 <= 'd0;
		in_data201 <= 'd0;
		in_data202 <= 'd0;
		in_data203 <= 'd0;
		in_data204 <= 'd0;
		in_data205 <= 'd0;
		in_data206 <= 'd0;
		in_data207 <= 'd0;
		in_data208 <= 'd0;
		in_data209 <= 'd0;
		in_data210 <= 'd0;
		in_data211 <= 'd0;
		in_data212 <= 'd0;
		in_data213 <= 'd0;
		in_data214 <= 'd0;
		in_data215 <= 'd0;
		in_data216 <= 'd0;
		in_data217 <= 'd0;
		in_data218 <= 'd0;
		in_data219 <= 'd0;
		in_data220 <= 'd0;
		in_data221 <= 'd0;
		in_data222 <= 'd0;
		in_data223 <= 'd0;
		in_data224 <= 'd0;
		in_data225 <= 'd0;
		in_data226 <= 'd0;
		in_data227 <= 'd0;
		in_data228 <= 'd0;
		in_data229 <= 'd0;
		in_data230 <= 'd0;
		in_data231 <= 'd0;
		in_data232 <= 'd0;
		in_data233 <= 'd0;
		in_data234 <= 'd0;
		in_data235 <= 'd0;
		in_data236 <= 'd0;
		in_data237 <= 'd0;
		in_data238 <= 'd0;
		in_data239 <= 'd0;
		in_data240 <= 'd0;
		in_data241 <= 'd0;
		in_data242 <= 'd0;
		in_data243 <= 'd0;
		in_data244 <= 'd0;
		in_data245 <= 'd0;
		in_data246 <= 'd0;
		in_data247 <= 'd0;
		in_data248 <= 'd0;
		in_data249 <= 'd0;
		in_data250 <= 'd0;
		in_data251 <= 'd0;
		in_data252 <= 'd0;
		in_data253 <= 'd0;
		in_data254 <= 'd0;
		in_data255 <= 'd0;
	end
	else begin
		if(in_valid) begin
			in_valid_flag <= 1'b1;
			input_index <= input_index + 'd1;
			IN_DATA(input_index) <= in_data;
		end
		else begin
			if(in_valid_flag) begin
				bubble_start_flag <= 1'b1;
			end
			else begin
				bubble_start_flag <= 1'b0;
			end
		end
	end
end



/*
 * Bubble Sort
 * -------------
 * - Break into ODD and EVEN parts
 * - INDEX of OUTER LOOP set to # of INPUTS (for now)
 */

reg				[7:0] outer_loop;
always @(posedge clk) begin
	if (!rst_n) begin
		outer_loop <= 'd0;		
	end
	else if (bubble_start_flag) begin
		if(outer_loop != input_index) begin
			outer_loop <= outer_loop + 1'b1;
		end
		else begin
			outer_loop <= outer_loop;
		end
	end
end


/*
 * Dump Output
 */
 reg			[7:0] output_index;
always @(posedge clk) begin
	if (!rst_n) begin
		output_index <= 'd0;		
	end
	else if (outer_loop == input_index) begin
		if (output_index < input_index) begin
			output_index <= output_index + 1'b1;
			out_data <= IN_DATA(output_index);
			out_valid <= 1'b1;
		end
		else begin
			out_data <= 'd0;
			out_valid <= 1'b0;
		end
	end
	else begin
		out_data <= 'd0;
		out_valid <= 1'b0;
	end
end



/*
 * Combinational Block for exchaging elements
 */

reg			[7:0] temp_even0;
reg			[7:0] temp_even1;
reg			[7:0] temp_even2;
reg			[7:0] temp_even3;
reg			[7:0] temp_even4;
reg			[7:0] temp_even5;
reg			[7:0] temp_even6;
reg			[7:0] temp_even7;
reg			[7:0] temp_even8;
reg			[7:0] temp_even9;
reg			[7:0] temp_even10;
reg			[7:0] temp_even11;
reg			[7:0] temp_even12;
reg			[7:0] temp_even13;
reg			[7:0] temp_even14;
reg			[7:0] temp_even15;
reg			[7:0] temp_even16;
reg			[7:0] temp_even17;
reg			[7:0] temp_even18;
reg			[7:0] temp_even19;
reg			[7:0] temp_even20;
reg			[7:0] temp_even21;
reg			[7:0] temp_even22;
reg			[7:0] temp_even23;
reg			[7:0] temp_even24;
reg			[7:0] temp_even25;
reg			[7:0] temp_even26;
reg			[7:0] temp_even27;
reg			[7:0] temp_even28;
reg			[7:0] temp_even29;
reg			[7:0] temp_even30;
reg			[7:0] temp_even31;
reg			[7:0] temp_even32;
reg			[7:0] temp_even33;
reg			[7:0] temp_even34;
reg			[7:0] temp_even35;
reg			[7:0] temp_even36;
reg			[7:0] temp_even37;
reg			[7:0] temp_even38;
reg			[7:0] temp_even39;
reg			[7:0] temp_even40;
reg			[7:0] temp_even41;
reg			[7:0] temp_even42;
reg			[7:0] temp_even43;
reg			[7:0] temp_even44;
reg			[7:0] temp_even45;
reg			[7:0] temp_even46;
reg			[7:0] temp_even47;
reg			[7:0] temp_even48;
reg			[7:0] temp_even49;
reg			[7:0] temp_even50;
reg			[7:0] temp_even51;
reg			[7:0] temp_even52;
reg			[7:0] temp_even53;
reg			[7:0] temp_even54;
reg			[7:0] temp_even55;
reg			[7:0] temp_even56;
reg			[7:0] temp_even57;
reg			[7:0] temp_even58;
reg			[7:0] temp_even59;
reg			[7:0] temp_even60;
reg			[7:0] temp_even61;
reg			[7:0] temp_even62;
reg			[7:0] temp_even63;
reg			[7:0] temp_even64;
reg			[7:0] temp_even65;
reg			[7:0] temp_even66;
reg			[7:0] temp_even67;
reg			[7:0] temp_even68;
reg			[7:0] temp_even69;
reg			[7:0] temp_even70;
reg			[7:0] temp_even71;
reg			[7:0] temp_even72;
reg			[7:0] temp_even73;
reg			[7:0] temp_even74;
reg			[7:0] temp_even75;
reg			[7:0] temp_even76;
reg			[7:0] temp_even77;
reg			[7:0] temp_even78;
reg			[7:0] temp_even79;
reg			[7:0] temp_even80;
reg			[7:0] temp_even81;
reg			[7:0] temp_even82;
reg			[7:0] temp_even83;
reg			[7:0] temp_even84;
reg			[7:0] temp_even85;
reg			[7:0] temp_even86;
reg			[7:0] temp_even87;
reg			[7:0] temp_even88;
reg			[7:0] temp_even89;
reg			[7:0] temp_even90;
reg			[7:0] temp_even91;
reg			[7:0] temp_even92;
reg			[7:0] temp_even93;
reg			[7:0] temp_even94;
reg			[7:0] temp_even95;
reg			[7:0] temp_even96;
reg			[7:0] temp_even97;
reg			[7:0] temp_even98;
reg			[7:0] temp_even99;
reg			[7:0] temp_even100;
reg			[7:0] temp_even101;
reg			[7:0] temp_even102;
reg			[7:0] temp_even103;
reg			[7:0] temp_even104;
reg			[7:0] temp_even105;
reg			[7:0] temp_even106;
reg			[7:0] temp_even107;
reg			[7:0] temp_even108;
reg			[7:0] temp_even109;
reg			[7:0] temp_even110;
reg			[7:0] temp_even111;
reg			[7:0] temp_even112;
reg			[7:0] temp_even113;
reg			[7:0] temp_even114;
reg			[7:0] temp_even115;
reg			[7:0] temp_even116;
reg			[7:0] temp_even117;
reg			[7:0] temp_even118;
reg			[7:0] temp_even119;
reg			[7:0] temp_even120;
reg			[7:0] temp_even121;
reg			[7:0] temp_even122;
reg			[7:0] temp_even123;
reg			[7:0] temp_even124;
reg			[7:0] temp_even125;
reg			[7:0] temp_even126;
reg			[7:0] temp_even127;
reg			[7:0] temp_even128;



reg			[7:0] temp_odd0;
reg			[7:0] temp_odd1;
reg			[7:0] temp_odd2;
reg			[7:0] temp_odd3;
reg			[7:0] temp_odd4;
reg			[7:0] temp_odd5;
reg			[7:0] temp_odd6;
reg			[7:0] temp_odd7;
reg			[7:0] temp_odd8;
reg			[7:0] temp_odd9;
reg			[7:0] temp_odd10;
reg			[7:0] temp_odd11;
reg			[7:0] temp_odd12;
reg			[7:0] temp_odd13;
reg			[7:0] temp_odd14;
reg			[7:0] temp_odd15;
reg			[7:0] temp_odd16;
reg			[7:0] temp_odd17;
reg			[7:0] temp_odd18;
reg			[7:0] temp_odd19;
reg			[7:0] temp_odd20;
reg			[7:0] temp_odd21;
reg			[7:0] temp_odd22;
reg			[7:0] temp_odd23;
reg			[7:0] temp_odd24;
reg			[7:0] temp_odd25;
reg			[7:0] temp_odd26;
reg			[7:0] temp_odd27;
reg			[7:0] temp_odd28;
reg			[7:0] temp_odd29;
reg			[7:0] temp_odd30;
reg			[7:0] temp_odd31;
reg			[7:0] temp_odd32;
reg			[7:0] temp_odd33;
reg			[7:0] temp_odd34;
reg			[7:0] temp_odd35;
reg			[7:0] temp_odd36;
reg			[7:0] temp_odd37;
reg			[7:0] temp_odd38;
reg			[7:0] temp_odd39;
reg			[7:0] temp_odd40;
reg			[7:0] temp_odd41;
reg			[7:0] temp_odd42;
reg			[7:0] temp_odd43;
reg			[7:0] temp_odd44;
reg			[7:0] temp_odd45;
reg			[7:0] temp_odd46;
reg			[7:0] temp_odd47;
reg			[7:0] temp_odd48;
reg			[7:0] temp_odd49;
reg			[7:0] temp_odd50;
reg			[7:0] temp_odd51;
reg			[7:0] temp_odd52;
reg			[7:0] temp_odd53;
reg			[7:0] temp_odd54;
reg			[7:0] temp_odd55;
reg			[7:0] temp_odd56;
reg			[7:0] temp_odd57;
reg			[7:0] temp_odd58;
reg			[7:0] temp_odd59;
reg			[7:0] temp_odd60;
reg			[7:0] temp_odd61;
reg			[7:0] temp_odd62;
reg			[7:0] temp_odd63;
reg			[7:0] temp_odd64;
reg			[7:0] temp_odd65;
reg			[7:0] temp_odd66;
reg			[7:0] temp_odd67;
reg			[7:0] temp_odd68;
reg			[7:0] temp_odd69;
reg			[7:0] temp_odd70;
reg			[7:0] temp_odd71;
reg			[7:0] temp_odd72;
reg			[7:0] temp_odd73;
reg			[7:0] temp_odd74;
reg			[7:0] temp_odd75;
reg			[7:0] temp_odd76;
reg			[7:0] temp_odd77;
reg			[7:0] temp_odd78;
reg			[7:0] temp_odd79;
reg			[7:0] temp_odd80;
reg			[7:0] temp_odd81;
reg			[7:0] temp_odd82;
reg			[7:0] temp_odd83;
reg			[7:0] temp_odd84;
reg			[7:0] temp_odd85;
reg			[7:0] temp_odd86;
reg			[7:0] temp_odd87;
reg			[7:0] temp_odd88;
reg			[7:0] temp_odd89;
reg			[7:0] temp_odd90;
reg			[7:0] temp_odd91;
reg			[7:0] temp_odd92;
reg			[7:0] temp_odd93;
reg			[7:0] temp_odd94;
reg			[7:0] temp_odd95;
reg			[7:0] temp_odd96;
reg			[7:0] temp_odd97;
reg			[7:0] temp_odd98;
reg			[7:0] temp_odd99;
reg			[7:0] temp_odd100;
reg			[7:0] temp_odd101;
reg			[7:0] temp_odd102;
reg			[7:0] temp_odd103;
reg			[7:0] temp_odd104;
reg			[7:0] temp_odd105;
reg			[7:0] temp_odd106;
reg			[7:0] temp_odd107;
reg			[7:0] temp_odd108;
reg			[7:0] temp_odd109;
reg			[7:0] temp_odd110;
reg			[7:0] temp_odd111;
reg			[7:0] temp_odd112;
reg			[7:0] temp_odd113;
reg			[7:0] temp_odd114;
reg			[7:0] temp_odd115;
reg			[7:0] temp_odd116;
reg			[7:0] temp_odd117;
reg			[7:0] temp_odd118;
reg			[7:0] temp_odd119;
reg			[7:0] temp_odd120;
reg			[7:0] temp_odd121;
reg			[7:0] temp_odd122;
reg			[7:0] temp_odd123;
reg			[7:0] temp_odd124;
reg			[7:0] temp_odd125;
reg			[7:0] temp_odd126;
reg			[7:0] temp_odd127;


/*
 * Swapping of Elements of Bubble Sort
 */

always @(*) begin
	if (bubble_start_flag) begin
		if(outer_loop[0:0] == 1'b1) begin //odd
			if(IN_DATA(1) < IN_DATA(2)) begin
				TEMP_ODD(1) = IN_DATA(1);
				IN_DATA(1) = IN_DATA(2);
				IN_DATA(2) = TEMP_ODD(1);
			end
			else begin
				TEMP_ODD(1) = 'd0;
			end
			if(IN_DATA(3) < IN_DATA(4)) begin
				TEMP_ODD(2) = IN_DATA(3);
				IN_DATA(3) = IN_DATA(4);
				IN_DATA(4) = TEMP_ODD(2);
			end
			else begin
				TEMP_ODD(2) = 'd0;
			end
			if(IN_DATA(5) < IN_DATA(6)) begin
				TEMP_ODD(3) = IN_DATA(5);
				IN_DATA(5) = IN_DATA(6);
				IN_DATA(6) = TEMP_ODD(3);
			end
			else begin
				TEMP_ODD(3) = 'd0;
			end
			if(IN_DATA(7) < IN_DATA(8)) begin
				TEMP_ODD(4) = IN_DATA(7);
				IN_DATA(7) = IN_DATA(8);
				IN_DATA(8) = TEMP_ODD(4);
			end
			else begin
				TEMP_ODD(4) = 'd0;
			end
			if(IN_DATA(9) < IN_DATA(10)) begin
				TEMP_ODD(5) = IN_DATA(9);
				IN_DATA(9) = IN_DATA(10);
				IN_DATA(10) = TEMP_ODD(5);
			end
			else begin
				TEMP_ODD(5) = 'd0;
			end
			if(IN_DATA(11) < IN_DATA(12)) begin
				TEMP_ODD(6) = IN_DATA(11);
				IN_DATA(11) = IN_DATA(12);
				IN_DATA(12) = TEMP_ODD(6);
			end
			else begin
				TEMP_ODD(6) = 'd0;
			end
			if(IN_DATA(13) < IN_DATA(14)) begin
				TEMP_ODD(7) = IN_DATA(13);
				IN_DATA(13) = IN_DATA(14);
				IN_DATA(14) = TEMP_ODD(7);
			end
			else begin
				TEMP_ODD(7) = 'd0;
			end
			if(IN_DATA(15) < IN_DATA(16)) begin
				TEMP_ODD(8) = IN_DATA(15);
				IN_DATA(15) = IN_DATA(16);
				IN_DATA(16) = TEMP_ODD(8);
			end
			else begin
				TEMP_ODD(8) = 'd0;
			end
			if(IN_DATA(17) < IN_DATA(18)) begin
				TEMP_ODD(9) = IN_DATA(17);
				IN_DATA(17) = IN_DATA(18);
				IN_DATA(18) = TEMP_ODD(9);
			end
			else begin
				TEMP_ODD(9) = 'd0;
			end
			if(IN_DATA(19) < IN_DATA(20)) begin
				TEMP_ODD(10) = IN_DATA(19);
				IN_DATA(19) = IN_DATA(20);
				IN_DATA(20) = TEMP_ODD(10);
			end
			else begin
				TEMP_ODD(10) = 'd0;
			end
			if(IN_DATA(21) < IN_DATA(22)) begin
				TEMP_ODD(11) = IN_DATA(21);
				IN_DATA(21) = IN_DATA(22);
				IN_DATA(22) = TEMP_ODD(11);
			end
			else begin
				TEMP_ODD(11) = 'd0;
			end
			if(IN_DATA(23) < IN_DATA(24)) begin
				TEMP_ODD(12) = IN_DATA(23);
				IN_DATA(23) = IN_DATA(24);
				IN_DATA(24) = TEMP_ODD(12);
			end
			else begin
				TEMP_ODD(12) = 'd0;
			end
			if(IN_DATA(25) < IN_DATA(26)) begin
				TEMP_ODD(13) = IN_DATA(25);
				IN_DATA(25) = IN_DATA(26);
				IN_DATA(26) = TEMP_ODD(13);
			end
			else begin
				TEMP_ODD(13) = 'd0;
			end
			if(IN_DATA(27) < IN_DATA(28)) begin
				TEMP_ODD(14) = IN_DATA(27);
				IN_DATA(27) = IN_DATA(28);
				IN_DATA(28) = TEMP_ODD(14);
			end
			else begin
				TEMP_ODD(14) = 'd0;
			end
			if(IN_DATA(29) < IN_DATA(30)) begin
				TEMP_ODD(15) = IN_DATA(29);
				IN_DATA(29) = IN_DATA(30);
				IN_DATA(30) = TEMP_ODD(15);
			end
			else begin
				TEMP_ODD(15) = 'd0;
			end
			if(IN_DATA(31) < IN_DATA(32)) begin
				TEMP_ODD(16) = IN_DATA(31);
				IN_DATA(31) = IN_DATA(32);
				IN_DATA(32) = TEMP_ODD(16);
			end
			else begin
				TEMP_ODD(16) = 'd0;
			end
			if(IN_DATA(33) < IN_DATA(34)) begin
				TEMP_ODD(17) = IN_DATA(33);
				IN_DATA(33) = IN_DATA(34);
				IN_DATA(34) = TEMP_ODD(17);
			end
			else begin
				TEMP_ODD(17) = 'd0;
			end
			if(IN_DATA(35) < IN_DATA(36)) begin
				TEMP_ODD(18) = IN_DATA(35);
				IN_DATA(35) = IN_DATA(36);
				IN_DATA(36) = TEMP_ODD(18);
			end
			else begin
				TEMP_ODD(18) = 'd0;
			end
			if(IN_DATA(37) < IN_DATA(38)) begin
				TEMP_ODD(19) = IN_DATA(37);
				IN_DATA(37) = IN_DATA(38);
				IN_DATA(38) = TEMP_ODD(19);
			end
			else begin
				TEMP_ODD(19) = 'd0;
			end
			if(IN_DATA(39) < IN_DATA(40)) begin
				TEMP_ODD(20) = IN_DATA(39);
				IN_DATA(39) = IN_DATA(40);
				IN_DATA(40) = TEMP_ODD(20);
			end
			else begin
				TEMP_ODD(20) = 'd0;
			end
			if(IN_DATA(41) < IN_DATA(42)) begin
				TEMP_ODD(21) = IN_DATA(41);
				IN_DATA(41) = IN_DATA(42);
				IN_DATA(42) = TEMP_ODD(21);
			end
			else begin
				TEMP_ODD(21) = 'd0;
			end
			if(IN_DATA(43) < IN_DATA(44)) begin
				TEMP_ODD(22) = IN_DATA(43);
				IN_DATA(43) = IN_DATA(44);
				IN_DATA(44) = TEMP_ODD(22);
			end
			else begin
				TEMP_ODD(22) = 'd0;
			end
			if(IN_DATA(45) < IN_DATA(46)) begin
				TEMP_ODD(23) = IN_DATA(45);
				IN_DATA(45) = IN_DATA(46);
				IN_DATA(46) = TEMP_ODD(23);
			end
			else begin
				TEMP_ODD(23) = 'd0;
			end
			if(IN_DATA(47) < IN_DATA(48)) begin
				TEMP_ODD(24) = IN_DATA(47);
				IN_DATA(47) = IN_DATA(48);
				IN_DATA(48) = TEMP_ODD(24);
			end
			else begin
				TEMP_ODD(24) = 'd0;
			end
			if(IN_DATA(49) < IN_DATA(50)) begin
				TEMP_ODD(25) = IN_DATA(49);
				IN_DATA(49) = IN_DATA(50);
				IN_DATA(50) = TEMP_ODD(25);
			end
			else begin
				TEMP_ODD(25) = 'd0;
			end
			if(IN_DATA(51) < IN_DATA(52)) begin
				TEMP_ODD(26) = IN_DATA(51);
				IN_DATA(51) = IN_DATA(52);
				IN_DATA(52) = TEMP_ODD(26);
			end
			else begin
				TEMP_ODD(26) = 'd0;
			end
			if(IN_DATA(53) < IN_DATA(54)) begin
				TEMP_ODD(27) = IN_DATA(53);
				IN_DATA(53) = IN_DATA(54);
				IN_DATA(54) = TEMP_ODD(27);
			end
			else begin
				TEMP_ODD(27) = 'd0;
			end
			if(IN_DATA(55) < IN_DATA(56)) begin
				TEMP_ODD(28) = IN_DATA(55);
				IN_DATA(55) = IN_DATA(56);
				IN_DATA(56) = TEMP_ODD(28);
			end
			else begin
				TEMP_ODD(28) = 'd0;
			end
			if(IN_DATA(57) < IN_DATA(58)) begin
				TEMP_ODD(29) = IN_DATA(57);
				IN_DATA(57) = IN_DATA(58);
				IN_DATA(58) = TEMP_ODD(29);
			end
			else begin
				TEMP_ODD(29) = 'd0;
			end
			if(IN_DATA(59) < IN_DATA(60)) begin
				TEMP_ODD(30) = IN_DATA(59);
				IN_DATA(59) = IN_DATA(60);
				IN_DATA(60) = TEMP_ODD(30);
			end
			else begin
				TEMP_ODD(30) = 'd0;
			end
			if(IN_DATA(61) < IN_DATA(62)) begin
				TEMP_ODD(31) = IN_DATA(61);
				IN_DATA(61) = IN_DATA(62);
				IN_DATA(62) = TEMP_ODD(31);
			end
			else begin
				TEMP_ODD(31) = 'd0;
			end
			if(IN_DATA(63) < IN_DATA(64)) begin
				TEMP_ODD(32) = IN_DATA(63);
				IN_DATA(63) = IN_DATA(64);
				IN_DATA(64) = TEMP_ODD(32);
			end
			else begin
				TEMP_ODD(32) = 'd0;
			end
			if(IN_DATA(65) < IN_DATA(66)) begin
				TEMP_ODD(33) = IN_DATA(65);
				IN_DATA(65) = IN_DATA(66);
				IN_DATA(66) = TEMP_ODD(33);
			end
			else begin
				TEMP_ODD(33) = 'd0;
			end
			if(IN_DATA(67) < IN_DATA(68)) begin
				TEMP_ODD(34) = IN_DATA(67);
				IN_DATA(67) = IN_DATA(68);
				IN_DATA(68) = TEMP_ODD(34);
			end
			else begin
				TEMP_ODD(34) = 'd0;
			end
			if(IN_DATA(69) < IN_DATA(70)) begin
				TEMP_ODD(35) = IN_DATA(69);
				IN_DATA(69) = IN_DATA(70);
				IN_DATA(70) = TEMP_ODD(35);
			end
			else begin
				TEMP_ODD(35) = 'd0;
			end
			if(IN_DATA(71) < IN_DATA(72)) begin
				TEMP_ODD(36) = IN_DATA(71);
				IN_DATA(71) = IN_DATA(72);
				IN_DATA(72) = TEMP_ODD(36);
			end
			else begin
				TEMP_ODD(36) = 'd0;
			end
			if(IN_DATA(73) < IN_DATA(74)) begin
				TEMP_ODD(37) = IN_DATA(73);
				IN_DATA(73) = IN_DATA(74);
				IN_DATA(74) = TEMP_ODD(37);
			end
			else begin
				TEMP_ODD(37) = 'd0;
			end
			if(IN_DATA(75) < IN_DATA(76)) begin
				TEMP_ODD(38) = IN_DATA(75);
				IN_DATA(75) = IN_DATA(76);
				IN_DATA(76) = TEMP_ODD(38);
			end
			else begin
				TEMP_ODD(38) = 'd0;
			end
			if(IN_DATA(77) < IN_DATA(78)) begin
				TEMP_ODD(39) = IN_DATA(77);
				IN_DATA(77) = IN_DATA(78);
				IN_DATA(78) = TEMP_ODD(39);
			end
			else begin
				TEMP_ODD(39) = 'd0;
			end
			if(IN_DATA(79) < IN_DATA(80)) begin
				TEMP_ODD(40) = IN_DATA(79);
				IN_DATA(79) = IN_DATA(80);
				IN_DATA(80) = TEMP_ODD(40);
			end
			else begin
				TEMP_ODD(40) = 'd0;
			end
			if(IN_DATA(81) < IN_DATA(82)) begin
				TEMP_ODD(41) = IN_DATA(81);
				IN_DATA(81) = IN_DATA(82);
				IN_DATA(82) = TEMP_ODD(41);
			end
			else begin
				TEMP_ODD(41) = 'd0;
			end
			if(IN_DATA(83) < IN_DATA(84)) begin
				TEMP_ODD(42) = IN_DATA(83);
				IN_DATA(83) = IN_DATA(84);
				IN_DATA(84) = TEMP_ODD(42);
			end
			else begin
				TEMP_ODD(42) = 'd0;
			end
			if(IN_DATA(85) < IN_DATA(86)) begin
				TEMP_ODD(43) = IN_DATA(85);
				IN_DATA(85) = IN_DATA(86);
				IN_DATA(86) = TEMP_ODD(43);
			end
			else begin
				TEMP_ODD(43) = 'd0;
			end
			if(IN_DATA(87) < IN_DATA(88)) begin
				TEMP_ODD(44) = IN_DATA(87);
				IN_DATA(87) = IN_DATA(88);
				IN_DATA(88) = TEMP_ODD(44);
			end
			else begin
				TEMP_ODD(44) = 'd0;
			end
			if(IN_DATA(89) < IN_DATA(90)) begin
				TEMP_ODD(45) = IN_DATA(89);
				IN_DATA(89) = IN_DATA(90);
				IN_DATA(90) = TEMP_ODD(45);
			end
			else begin
				TEMP_ODD(45) = 'd0;
			end
			if(IN_DATA(91) < IN_DATA(92)) begin
				TEMP_ODD(46) = IN_DATA(91);
				IN_DATA(91) = IN_DATA(92);
				IN_DATA(92) = TEMP_ODD(46);
			end
			else begin
				TEMP_ODD(46) = 'd0;
			end
			if(IN_DATA(93) < IN_DATA(94)) begin
				TEMP_ODD(47) = IN_DATA(93);
				IN_DATA(93) = IN_DATA(94);
				IN_DATA(94) = TEMP_ODD(47);
			end
			else begin
				TEMP_ODD(47) = 'd0;
			end
			if(IN_DATA(95) < IN_DATA(96)) begin
				TEMP_ODD(48) = IN_DATA(95);
				IN_DATA(95) = IN_DATA(96);
				IN_DATA(96) = TEMP_ODD(48);
			end
			else begin
				TEMP_ODD(48) = 'd0;
			end
			if(IN_DATA(97) < IN_DATA(98)) begin
				TEMP_ODD(49) = IN_DATA(97);
				IN_DATA(97) = IN_DATA(98);
				IN_DATA(98) = TEMP_ODD(49);
			end
			else begin
				TEMP_ODD(49) = 'd0;
			end
			if(IN_DATA(99) < IN_DATA(100)) begin
				TEMP_ODD(50) = IN_DATA(99);
				IN_DATA(99) = IN_DATA(100);
				IN_DATA(100) = TEMP_ODD(50);
			end
			else begin
				TEMP_ODD(50) = 'd0;
			end
			if(IN_DATA(101) < IN_DATA(102)) begin
				TEMP_ODD(51) = IN_DATA(101);
				IN_DATA(101) = IN_DATA(102);
				IN_DATA(102) = TEMP_ODD(51);
			end
			else begin
				TEMP_ODD(51) = 'd0;
			end
			if(IN_DATA(103) < IN_DATA(104)) begin
				TEMP_ODD(52) = IN_DATA(103);
				IN_DATA(103) = IN_DATA(104);
				IN_DATA(104) = TEMP_ODD(52);
			end
			else begin
				TEMP_ODD(52) = 'd0;
			end
			if(IN_DATA(105) < IN_DATA(106)) begin
				TEMP_ODD(53) = IN_DATA(105);
				IN_DATA(105) = IN_DATA(106);
				IN_DATA(106) = TEMP_ODD(53);
			end
			else begin
				TEMP_ODD(53) = 'd0;
			end
			if(IN_DATA(107) < IN_DATA(108)) begin
				TEMP_ODD(54) = IN_DATA(107);
				IN_DATA(107) = IN_DATA(108);
				IN_DATA(108) = TEMP_ODD(54);
			end
			else begin
				TEMP_ODD(54) = 'd0;
			end
			if(IN_DATA(109) < IN_DATA(110)) begin
				TEMP_ODD(55) = IN_DATA(109);
				IN_DATA(109) = IN_DATA(110);
				IN_DATA(110) = TEMP_ODD(55);
			end
			else begin
				TEMP_ODD(55) = 'd0;
			end
			if(IN_DATA(111) < IN_DATA(112)) begin
				TEMP_ODD(56) = IN_DATA(111);
				IN_DATA(111) = IN_DATA(112);
				IN_DATA(112) = TEMP_ODD(56);
			end
			else begin
				TEMP_ODD(56) = 'd0;
			end
			if(IN_DATA(113) < IN_DATA(114)) begin
				TEMP_ODD(57) = IN_DATA(113);
				IN_DATA(113) = IN_DATA(114);
				IN_DATA(114) = TEMP_ODD(57);
			end
			else begin
				TEMP_ODD(57) = 'd0;
			end
			if(IN_DATA(115) < IN_DATA(116)) begin
				TEMP_ODD(58) = IN_DATA(115);
				IN_DATA(115) = IN_DATA(116);
				IN_DATA(116) = TEMP_ODD(58);
			end
			else begin
				TEMP_ODD(58) = 'd0;
			end
			if(IN_DATA(117) < IN_DATA(118)) begin
				TEMP_ODD(59) = IN_DATA(117);
				IN_DATA(117) = IN_DATA(118);
				IN_DATA(118) = TEMP_ODD(59);
			end
			else begin
				TEMP_ODD(59) = 'd0;
			end
			if(IN_DATA(119) < IN_DATA(120)) begin
				TEMP_ODD(60) = IN_DATA(119);
				IN_DATA(119) = IN_DATA(120);
				IN_DATA(120) = TEMP_ODD(60);
			end
			else begin
				TEMP_ODD(60) = 'd0;
			end
			if(IN_DATA(121) < IN_DATA(122)) begin
				TEMP_ODD(61) = IN_DATA(121);
				IN_DATA(121) = IN_DATA(122);
				IN_DATA(122) = TEMP_ODD(61);
			end
			else begin
				TEMP_ODD(61) = 'd0;
			end
			if(IN_DATA(123) < IN_DATA(124)) begin
				TEMP_ODD(62) = IN_DATA(123);
				IN_DATA(123) = IN_DATA(124);
				IN_DATA(124) = TEMP_ODD(62);
			end
			else begin
				TEMP_ODD(62) = 'd0;
			end
			if(IN_DATA(125) < IN_DATA(126)) begin
				TEMP_ODD(63) = IN_DATA(125);
				IN_DATA(125) = IN_DATA(126);
				IN_DATA(126) = TEMP_ODD(63);
			end
			else begin
				TEMP_ODD(63) = 'd0;
			end
			if(IN_DATA(127) < IN_DATA(128)) begin
				TEMP_ODD(64) = IN_DATA(127);
				IN_DATA(127) = IN_DATA(128);
				IN_DATA(128) = TEMP_ODD(64);
			end
			else begin
				TEMP_ODD(64) = 'd0;
			end
			if(IN_DATA(129) < IN_DATA(130)) begin
				TEMP_ODD(65) = IN_DATA(129);
				IN_DATA(129) = IN_DATA(130);
				IN_DATA(130) = TEMP_ODD(65);
			end
			else begin
				TEMP_ODD(65) = 'd0;
			end
			if(IN_DATA(131) < IN_DATA(132)) begin
				TEMP_ODD(66) = IN_DATA(131);
				IN_DATA(131) = IN_DATA(132);
				IN_DATA(132) = TEMP_ODD(66);
			end
			else begin
				TEMP_ODD(66) = 'd0;
			end
			if(IN_DATA(133) < IN_DATA(134)) begin
				TEMP_ODD(67) = IN_DATA(133);
				IN_DATA(133) = IN_DATA(134);
				IN_DATA(134) = TEMP_ODD(67);
			end
			else begin
				TEMP_ODD(67) = 'd0;
			end
			if(IN_DATA(135) < IN_DATA(136)) begin
				TEMP_ODD(68) = IN_DATA(135);
				IN_DATA(135) = IN_DATA(136);
				IN_DATA(136) = TEMP_ODD(68);
			end
			else begin
				TEMP_ODD(68) = 'd0;
			end
			if(IN_DATA(137) < IN_DATA(138)) begin
				TEMP_ODD(69) = IN_DATA(137);
				IN_DATA(137) = IN_DATA(138);
				IN_DATA(138) = TEMP_ODD(69);
			end
			else begin
				TEMP_ODD(69) = 'd0;
			end
			if(IN_DATA(139) < IN_DATA(140)) begin
				TEMP_ODD(70) = IN_DATA(139);
				IN_DATA(139) = IN_DATA(140);
				IN_DATA(140) = TEMP_ODD(70);
			end
			else begin
				TEMP_ODD(70) = 'd0;
			end
			if(IN_DATA(141) < IN_DATA(142)) begin
				TEMP_ODD(71) = IN_DATA(141);
				IN_DATA(141) = IN_DATA(142);
				IN_DATA(142) = TEMP_ODD(71);
			end
			else begin
				TEMP_ODD(71) = 'd0;
			end
			if(IN_DATA(143) < IN_DATA(144)) begin
				TEMP_ODD(72) = IN_DATA(143);
				IN_DATA(143) = IN_DATA(144);
				IN_DATA(144) = TEMP_ODD(72);
			end
			else begin
				TEMP_ODD(72) = 'd0;
			end
			if(IN_DATA(145) < IN_DATA(146)) begin
				TEMP_ODD(73) = IN_DATA(145);
				IN_DATA(145) = IN_DATA(146);
				IN_DATA(146) = TEMP_ODD(73);
			end
			else begin
				TEMP_ODD(73) = 'd0;
			end
			if(IN_DATA(147) < IN_DATA(148)) begin
				TEMP_ODD(74) = IN_DATA(147);
				IN_DATA(147) = IN_DATA(148);
				IN_DATA(148) = TEMP_ODD(74);
			end
			else begin
				TEMP_ODD(74) = 'd0;
			end
			if(IN_DATA(149) < IN_DATA(150)) begin
				TEMP_ODD(75) = IN_DATA(149);
				IN_DATA(149) = IN_DATA(150);
				IN_DATA(150) = TEMP_ODD(75);
			end
			else begin
				TEMP_ODD(75) = 'd0;
			end
			if(IN_DATA(151) < IN_DATA(152)) begin
				TEMP_ODD(76) = IN_DATA(151);
				IN_DATA(151) = IN_DATA(152);
				IN_DATA(152) = TEMP_ODD(76);
			end
			else begin
				TEMP_ODD(76) = 'd0;
			end
			if(IN_DATA(153) < IN_DATA(154)) begin
				TEMP_ODD(77) = IN_DATA(153);
				IN_DATA(153) = IN_DATA(154);
				IN_DATA(154) = TEMP_ODD(77);
			end
			else begin
				TEMP_ODD(77) = 'd0;
			end
			if(IN_DATA(155) < IN_DATA(156)) begin
				TEMP_ODD(78) = IN_DATA(155);
				IN_DATA(155) = IN_DATA(156);
				IN_DATA(156) = TEMP_ODD(78);
			end
			else begin
				TEMP_ODD(78) = 'd0;
			end
			if(IN_DATA(157) < IN_DATA(158)) begin
				TEMP_ODD(79) = IN_DATA(157);
				IN_DATA(157) = IN_DATA(158);
				IN_DATA(158) = TEMP_ODD(79);
			end
			else begin
				TEMP_ODD(79) = 'd0;
			end
			if(IN_DATA(159) < IN_DATA(160)) begin
				TEMP_ODD(80) = IN_DATA(159);
				IN_DATA(159) = IN_DATA(160);
				IN_DATA(160) = TEMP_ODD(80);
			end
			else begin
				TEMP_ODD(80) = 'd0;
			end
			if(IN_DATA(161) < IN_DATA(162)) begin
				TEMP_ODD(81) = IN_DATA(161);
				IN_DATA(161) = IN_DATA(162);
				IN_DATA(162) = TEMP_ODD(81);
			end
			else begin
				TEMP_ODD(81) = 'd0;
			end
			if(IN_DATA(163) < IN_DATA(164)) begin
				TEMP_ODD(82) = IN_DATA(163);
				IN_DATA(163) = IN_DATA(164);
				IN_DATA(164) = TEMP_ODD(82);
			end
			else begin
				TEMP_ODD(82) = 'd0;
			end
			if(IN_DATA(165) < IN_DATA(166)) begin
				TEMP_ODD(83) = IN_DATA(165);
				IN_DATA(165) = IN_DATA(166);
				IN_DATA(166) = TEMP_ODD(83);
			end
			else begin
				TEMP_ODD(83) = 'd0;
			end
			if(IN_DATA(167) < IN_DATA(168)) begin
				TEMP_ODD(84) = IN_DATA(167);
				IN_DATA(167) = IN_DATA(168);
				IN_DATA(168) = TEMP_ODD(84);
			end
			else begin
				TEMP_ODD(84) = 'd0;
			end
			if(IN_DATA(169) < IN_DATA(170)) begin
				TEMP_ODD(85) = IN_DATA(169);
				IN_DATA(169) = IN_DATA(170);
				IN_DATA(170) = TEMP_ODD(85);
			end
			else begin
				TEMP_ODD(85) = 'd0;
			end
			if(IN_DATA(171) < IN_DATA(172)) begin
				TEMP_ODD(86) = IN_DATA(171);
				IN_DATA(171) = IN_DATA(172);
				IN_DATA(172) = TEMP_ODD(86);
			end
			else begin
				TEMP_ODD(86) = 'd0;
			end
			if(IN_DATA(173) < IN_DATA(174)) begin
				TEMP_ODD(87) = IN_DATA(173);
				IN_DATA(173) = IN_DATA(174);
				IN_DATA(174) = TEMP_ODD(87);
			end
			else begin
				TEMP_ODD(87) = 'd0;
			end
			if(IN_DATA(175) < IN_DATA(176)) begin
				TEMP_ODD(88) = IN_DATA(175);
				IN_DATA(175) = IN_DATA(176);
				IN_DATA(176) = TEMP_ODD(88);
			end
			else begin
				TEMP_ODD(88) = 'd0;
			end
			if(IN_DATA(177) < IN_DATA(178)) begin
				TEMP_ODD(89) = IN_DATA(177);
				IN_DATA(177) = IN_DATA(178);
				IN_DATA(178) = TEMP_ODD(89);
			end
			else begin
				TEMP_ODD(89) = 'd0;
			end
			if(IN_DATA(179) < IN_DATA(180)) begin
				TEMP_ODD(90) = IN_DATA(179);
				IN_DATA(179) = IN_DATA(180);
				IN_DATA(180) = TEMP_ODD(90);
			end
			else begin
				TEMP_ODD(90) = 'd0;
			end
			if(IN_DATA(181) < IN_DATA(182)) begin
				TEMP_ODD(91) = IN_DATA(181);
				IN_DATA(181) = IN_DATA(182);
				IN_DATA(182) = TEMP_ODD(91);
			end
			else begin
				TEMP_ODD(91) = 'd0;
			end
			if(IN_DATA(183) < IN_DATA(184)) begin
				TEMP_ODD(92) = IN_DATA(183);
				IN_DATA(183) = IN_DATA(184);
				IN_DATA(184) = TEMP_ODD(92);
			end
			else begin
				TEMP_ODD(92) = 'd0;
			end
			if(IN_DATA(185) < IN_DATA(186)) begin
				TEMP_ODD(93) = IN_DATA(185);
				IN_DATA(185) = IN_DATA(186);
				IN_DATA(186) = TEMP_ODD(93);
			end
			else begin
				TEMP_ODD(93) = 'd0;
			end
			if(IN_DATA(187) < IN_DATA(188)) begin
				TEMP_ODD(94) = IN_DATA(187);
				IN_DATA(187) = IN_DATA(188);
				IN_DATA(188) = TEMP_ODD(94);
			end
			else begin
				TEMP_ODD(94) = 'd0;
			end
			if(IN_DATA(189) < IN_DATA(190)) begin
				TEMP_ODD(95) = IN_DATA(189);
				IN_DATA(189) = IN_DATA(190);
				IN_DATA(190) = TEMP_ODD(95);
			end
			else begin
				TEMP_ODD(95) = 'd0;
			end
			if(IN_DATA(191) < IN_DATA(192)) begin
				TEMP_ODD(96) = IN_DATA(191);
				IN_DATA(191) = IN_DATA(192);
				IN_DATA(192) = TEMP_ODD(96);
			end
			else begin
				TEMP_ODD(96) = 'd0;
			end
			if(IN_DATA(193) < IN_DATA(194)) begin
				TEMP_ODD(97) = IN_DATA(193);
				IN_DATA(193) = IN_DATA(194);
				IN_DATA(194) = TEMP_ODD(97);
			end
			else begin
				TEMP_ODD(97) = 'd0;
			end
			if(IN_DATA(195) < IN_DATA(196)) begin
				TEMP_ODD(98) = IN_DATA(195);
				IN_DATA(195) = IN_DATA(196);
				IN_DATA(196) = TEMP_ODD(98);
			end
			else begin
				TEMP_ODD(98) = 'd0;
			end
			if(IN_DATA(197) < IN_DATA(198)) begin
				TEMP_ODD(99) = IN_DATA(197);
				IN_DATA(197) = IN_DATA(198);
				IN_DATA(198) = TEMP_ODD(99);
			end
			else begin
				TEMP_ODD(99) = 'd0;
			end
			if(IN_DATA(199) < IN_DATA(200)) begin
				TEMP_ODD(100) = IN_DATA(199);
				IN_DATA(199) = IN_DATA(200);
				IN_DATA(200) = TEMP_ODD(100);
			end
			else begin
				TEMP_ODD(100) = 'd0;
			end
			if(IN_DATA(201) < IN_DATA(202)) begin
				TEMP_ODD(101) = IN_DATA(201);
				IN_DATA(201) = IN_DATA(202);
				IN_DATA(202) = TEMP_ODD(101);
			end
			else begin
				TEMP_ODD(101) = 'd0;
			end
			if(IN_DATA(203) < IN_DATA(204)) begin
				TEMP_ODD(102) = IN_DATA(203);
				IN_DATA(203) = IN_DATA(204);
				IN_DATA(204) = TEMP_ODD(102);
			end
			else begin
				TEMP_ODD(102) = 'd0;
			end
			if(IN_DATA(205) < IN_DATA(206)) begin
				TEMP_ODD(103) = IN_DATA(205);
				IN_DATA(205) = IN_DATA(206);
				IN_DATA(206) = TEMP_ODD(103);
			end
			else begin
				TEMP_ODD(103) = 'd0;
			end
			if(IN_DATA(207) < IN_DATA(208)) begin
				TEMP_ODD(104) = IN_DATA(207);
				IN_DATA(207) = IN_DATA(208);
				IN_DATA(208) = TEMP_ODD(104);
			end
			else begin
				TEMP_ODD(104) = 'd0;
			end
			if(IN_DATA(209) < IN_DATA(210)) begin
				TEMP_ODD(105) = IN_DATA(209);
				IN_DATA(209) = IN_DATA(210);
				IN_DATA(210) = TEMP_ODD(105);
			end
			else begin
				TEMP_ODD(105) = 'd0;
			end
			if(IN_DATA(211) < IN_DATA(212)) begin
				TEMP_ODD(106) = IN_DATA(211);
				IN_DATA(211) = IN_DATA(212);
				IN_DATA(212) = TEMP_ODD(106);
			end
			else begin
				TEMP_ODD(106) = 'd0;
			end
			if(IN_DATA(213) < IN_DATA(214)) begin
				TEMP_ODD(107) = IN_DATA(213);
				IN_DATA(213) = IN_DATA(214);
				IN_DATA(214) = TEMP_ODD(107);
			end
			else begin
				TEMP_ODD(107) = 'd0;
			end
			if(IN_DATA(215) < IN_DATA(216)) begin
				TEMP_ODD(108) = IN_DATA(215);
				IN_DATA(215) = IN_DATA(216);
				IN_DATA(216) = TEMP_ODD(108);
			end
			else begin
				TEMP_ODD(108) = 'd0;
			end
			if(IN_DATA(217) < IN_DATA(218)) begin
				TEMP_ODD(109) = IN_DATA(217);
				IN_DATA(217) = IN_DATA(218);
				IN_DATA(218) = TEMP_ODD(109);
			end
			else begin
				TEMP_ODD(109) = 'd0;
			end
			if(IN_DATA(219) < IN_DATA(220)) begin
				TEMP_ODD(110) = IN_DATA(219);
				IN_DATA(219) = IN_DATA(220);
				IN_DATA(220) = TEMP_ODD(110);
			end
			else begin
				TEMP_ODD(110) = 'd0;
			end
			if(IN_DATA(221) < IN_DATA(222)) begin
				TEMP_ODD(111) = IN_DATA(221);
				IN_DATA(221) = IN_DATA(222);
				IN_DATA(222) = TEMP_ODD(111);
			end
			else begin
				TEMP_ODD(111) = 'd0;
			end
			if(IN_DATA(223) < IN_DATA(224)) begin
				TEMP_ODD(112) = IN_DATA(223);
				IN_DATA(223) = IN_DATA(224);
				IN_DATA(224) = TEMP_ODD(112);
			end
			else begin
				TEMP_ODD(112) = 'd0;
			end
			if(IN_DATA(225) < IN_DATA(226)) begin
				TEMP_ODD(113) = IN_DATA(225);
				IN_DATA(225) = IN_DATA(226);
				IN_DATA(226) = TEMP_ODD(113);
			end
			else begin
				TEMP_ODD(113) = 'd0;
			end
			if(IN_DATA(227) < IN_DATA(228)) begin
				TEMP_ODD(114) = IN_DATA(227);
				IN_DATA(227) = IN_DATA(228);
				IN_DATA(228) = TEMP_ODD(114);
			end
			else begin
				TEMP_ODD(114) = 'd0;
			end
			if(IN_DATA(229) < IN_DATA(230)) begin
				TEMP_ODD(115) = IN_DATA(229);
				IN_DATA(229) = IN_DATA(230);
				IN_DATA(230) = TEMP_ODD(115);
			end
			else begin
				TEMP_ODD(115) = 'd0;
			end
			if(IN_DATA(231) < IN_DATA(232)) begin
				TEMP_ODD(116) = IN_DATA(231);
				IN_DATA(231) = IN_DATA(232);
				IN_DATA(232) = TEMP_ODD(116);
			end
			else begin
				TEMP_ODD(116) = 'd0;
			end
			if(IN_DATA(233) < IN_DATA(234)) begin
				TEMP_ODD(117) = IN_DATA(233);
				IN_DATA(233) = IN_DATA(234);
				IN_DATA(234) = TEMP_ODD(117);
			end
			else begin
				TEMP_ODD(117) = 'd0;
			end
			if(IN_DATA(235) < IN_DATA(236)) begin
				TEMP_ODD(118) = IN_DATA(235);
				IN_DATA(235) = IN_DATA(236);
				IN_DATA(236) = TEMP_ODD(118);
			end
			else begin
				TEMP_ODD(118) = 'd0;
			end
			if(IN_DATA(237) < IN_DATA(238)) begin
				TEMP_ODD(119) = IN_DATA(237);
				IN_DATA(237) = IN_DATA(238);
				IN_DATA(238) = TEMP_ODD(119);
			end
			else begin
				TEMP_ODD(119) = 'd0;
			end
			if(IN_DATA(239) < IN_DATA(240)) begin
				TEMP_ODD(120) = IN_DATA(239);
				IN_DATA(239) = IN_DATA(240);
				IN_DATA(240) = TEMP_ODD(120);
			end
			else begin
				TEMP_ODD(120) = 'd0;
			end
			if(IN_DATA(241) < IN_DATA(242)) begin
				TEMP_ODD(121) = IN_DATA(241);
				IN_DATA(241) = IN_DATA(242);
				IN_DATA(242) = TEMP_ODD(121);
			end
			else begin
				TEMP_ODD(121) = 'd0;
			end
			if(IN_DATA(243) < IN_DATA(244)) begin
				TEMP_ODD(122) = IN_DATA(243);
				IN_DATA(243) = IN_DATA(244);
				IN_DATA(244) = TEMP_ODD(122);
			end
			else begin
				TEMP_ODD(122) = 'd0;
			end
			if(IN_DATA(245) < IN_DATA(246)) begin
				TEMP_ODD(123) = IN_DATA(245);
				IN_DATA(245) = IN_DATA(246);
				IN_DATA(246) = TEMP_ODD(123);
			end
			else begin
				TEMP_ODD(123) = 'd0;
			end
			if(IN_DATA(247) < IN_DATA(248)) begin
				TEMP_ODD(124) = IN_DATA(247);
				IN_DATA(247) = IN_DATA(248);
				IN_DATA(248) = TEMP_ODD(124);
			end
			else begin
				TEMP_ODD(124) = 'd0;
			end
			if(IN_DATA(249) < IN_DATA(250)) begin
				TEMP_ODD(125) = IN_DATA(249);
				IN_DATA(249) = IN_DATA(250);
				IN_DATA(250) = TEMP_ODD(125);
			end
			else begin
				TEMP_ODD(125) = 'd0;
			end
			if(IN_DATA(251) < IN_DATA(252)) begin
				TEMP_ODD(126) = IN_DATA(251);
				IN_DATA(251) = IN_DATA(252);
				IN_DATA(252) = TEMP_ODD(126);
			end
			else begin
				TEMP_ODD(126) = 'd0;
			end
			if(IN_DATA(253) < IN_DATA(254)) begin
				TEMP_ODD(127) = IN_DATA(253);
				IN_DATA(253) = IN_DATA(254);
				IN_DATA(254) = TEMP_ODD(127);
			end
			else begin
				TEMP_ODD(127) = 'd0;
			end
		end
		else begin //even
			if(IN_DATA(0) < IN_DATA(1)) begin
				TEMP_EVEN(1) = IN_DATA(0);
				IN_DATA(0) = IN_DATA(1);
				IN_DATA(1) = TEMP_EVEN(1);
			end
			else begin
				TEMP_EVEN(1) = 'd0;
			end
			if(IN_DATA(2) < IN_DATA(3)) begin
				TEMP_EVEN(2) = IN_DATA(2);
				IN_DATA(2) = IN_DATA(3);
				IN_DATA(3) = TEMP_EVEN(2);
			end
			else begin
				TEMP_EVEN(2) = 'd0;
			end
			if(IN_DATA(4) < IN_DATA(5)) begin
				TEMP_EVEN(3) = IN_DATA(4);
				IN_DATA(4) = IN_DATA(5);
				IN_DATA(5) = TEMP_EVEN(3);
			end
			else begin
				TEMP_EVEN(3) = 'd0;
			end
			if(IN_DATA(6) < IN_DATA(7)) begin
				TEMP_EVEN(4) = IN_DATA(6);
				IN_DATA(6) = IN_DATA(7);
				IN_DATA(7) = TEMP_EVEN(4);
			end
			else begin
				TEMP_EVEN(4) = 'd0;
			end
			if(IN_DATA(8) < IN_DATA(9)) begin
				TEMP_EVEN(5) = IN_DATA(8);
				IN_DATA(8) = IN_DATA(9);
				IN_DATA(9) = TEMP_EVEN(5);
			end
			else begin
				TEMP_EVEN(5) = 'd0;
			end
			if(IN_DATA(10) < IN_DATA(11)) begin
				TEMP_EVEN(6) = IN_DATA(10);
				IN_DATA(10) = IN_DATA(11);
				IN_DATA(11) = TEMP_EVEN(6);
			end
			else begin
				TEMP_EVEN(6) = 'd0;
			end
			if(IN_DATA(12) < IN_DATA(13)) begin
				TEMP_EVEN(7) = IN_DATA(12);
				IN_DATA(12) = IN_DATA(13);
				IN_DATA(13) = TEMP_EVEN(7);
			end
			else begin
				TEMP_EVEN(7) = 'd0;
			end
			if(IN_DATA(14) < IN_DATA(15)) begin
				TEMP_EVEN(8) = IN_DATA(14);
				IN_DATA(14) = IN_DATA(15);
				IN_DATA(15) = TEMP_EVEN(8);
			end
			else begin
				TEMP_EVEN(8) = 'd0;
			end
			if(IN_DATA(16) < IN_DATA(17)) begin
				TEMP_EVEN(9) = IN_DATA(16);
				IN_DATA(16) = IN_DATA(17);
				IN_DATA(17) = TEMP_EVEN(9);
			end
			else begin
				TEMP_EVEN(9) = 'd0;
			end
			if(IN_DATA(18) < IN_DATA(19)) begin
				TEMP_EVEN(10) = IN_DATA(18);
				IN_DATA(18) = IN_DATA(19);
				IN_DATA(19) = TEMP_EVEN(10);
			end
			else begin
				TEMP_EVEN(10) = 'd0;
			end
			if(IN_DATA(20) < IN_DATA(21)) begin
				TEMP_EVEN(11) = IN_DATA(20);
				IN_DATA(20) = IN_DATA(21);
				IN_DATA(21) = TEMP_EVEN(11);
			end
			else begin
				TEMP_EVEN(11) = 'd0;
			end
			if(IN_DATA(22) < IN_DATA(23)) begin
				TEMP_EVEN(12) = IN_DATA(22);
				IN_DATA(22) = IN_DATA(23);
				IN_DATA(23) = TEMP_EVEN(12);
			end
			else begin
				TEMP_EVEN(12) = 'd0;
			end
			if(IN_DATA(24) < IN_DATA(25)) begin
				TEMP_EVEN(13) = IN_DATA(24);
				IN_DATA(24) = IN_DATA(25);
				IN_DATA(25) = TEMP_EVEN(13);
			end
			else begin
				TEMP_EVEN(13) = 'd0;
			end
			if(IN_DATA(26) < IN_DATA(27)) begin
				TEMP_EVEN(14) = IN_DATA(26);
				IN_DATA(26) = IN_DATA(27);
				IN_DATA(27) = TEMP_EVEN(14);
			end
			else begin
				TEMP_EVEN(14) = 'd0;
			end
			if(IN_DATA(28) < IN_DATA(29)) begin
				TEMP_EVEN(15) = IN_DATA(28);
				IN_DATA(28) = IN_DATA(29);
				IN_DATA(29) = TEMP_EVEN(15);
			end
			else begin
				TEMP_EVEN(15) = 'd0;
			end
			if(IN_DATA(30) < IN_DATA(31)) begin
				TEMP_EVEN(16) = IN_DATA(30);
				IN_DATA(30) = IN_DATA(31);
				IN_DATA(31) = TEMP_EVEN(16);
			end
			else begin
				TEMP_EVEN(16) = 'd0;
			end
			if(IN_DATA(32) < IN_DATA(33)) begin
				TEMP_EVEN(17) = IN_DATA(32);
				IN_DATA(32) = IN_DATA(33);
				IN_DATA(33) = TEMP_EVEN(17);
			end
			else begin
				TEMP_EVEN(17) = 'd0;
			end
			if(IN_DATA(34) < IN_DATA(35)) begin
				TEMP_EVEN(18) = IN_DATA(34);
				IN_DATA(34) = IN_DATA(35);
				IN_DATA(35) = TEMP_EVEN(18);
			end
			else begin
				TEMP_EVEN(18) = 'd0;
			end
			if(IN_DATA(36) < IN_DATA(37)) begin
				TEMP_EVEN(19) = IN_DATA(36);
				IN_DATA(36) = IN_DATA(37);
				IN_DATA(37) = TEMP_EVEN(19);
			end
			else begin
				TEMP_EVEN(19) = 'd0;
			end
			if(IN_DATA(38) < IN_DATA(39)) begin
				TEMP_EVEN(20) = IN_DATA(38);
				IN_DATA(38) = IN_DATA(39);
				IN_DATA(39) = TEMP_EVEN(20);
			end
			else begin
				TEMP_EVEN(20) = 'd0;
			end
			if(IN_DATA(40) < IN_DATA(41)) begin
				TEMP_EVEN(21) = IN_DATA(40);
				IN_DATA(40) = IN_DATA(41);
				IN_DATA(41) = TEMP_EVEN(21);
			end
			else begin
				TEMP_EVEN(21) = 'd0;
			end
			if(IN_DATA(42) < IN_DATA(43)) begin
				TEMP_EVEN(22) = IN_DATA(42);
				IN_DATA(42) = IN_DATA(43);
				IN_DATA(43) = TEMP_EVEN(22);
			end
			else begin
				TEMP_EVEN(22) = 'd0;
			end
			if(IN_DATA(44) < IN_DATA(45)) begin
				TEMP_EVEN(23) = IN_DATA(44);
				IN_DATA(44) = IN_DATA(45);
				IN_DATA(45) = TEMP_EVEN(23);
			end
			else begin
				TEMP_EVEN(23) = 'd0;
			end
			if(IN_DATA(46) < IN_DATA(47)) begin
				TEMP_EVEN(24) = IN_DATA(46);
				IN_DATA(46) = IN_DATA(47);
				IN_DATA(47) = TEMP_EVEN(24);
			end
			else begin
				TEMP_EVEN(24) = 'd0;
			end
			if(IN_DATA(48) < IN_DATA(49)) begin
				TEMP_EVEN(25) = IN_DATA(48);
				IN_DATA(48) = IN_DATA(49);
				IN_DATA(49) = TEMP_EVEN(25);
			end
			else begin
				TEMP_EVEN(25) = 'd0;
			end
			if(IN_DATA(50) < IN_DATA(51)) begin
				TEMP_EVEN(26) = IN_DATA(50);
				IN_DATA(50) = IN_DATA(51);
				IN_DATA(51) = TEMP_EVEN(26);
			end
			else begin
				TEMP_EVEN(26) = 'd0;
			end
			if(IN_DATA(52) < IN_DATA(53)) begin
				TEMP_EVEN(27) = IN_DATA(52);
				IN_DATA(52) = IN_DATA(53);
				IN_DATA(53) = TEMP_EVEN(27);
			end
			else begin
				TEMP_EVEN(27) = 'd0;
			end
			if(IN_DATA(54) < IN_DATA(55)) begin
				TEMP_EVEN(28) = IN_DATA(54);
				IN_DATA(54) = IN_DATA(55);
				IN_DATA(55) = TEMP_EVEN(28);
			end
			else begin
				TEMP_EVEN(28) = 'd0;
			end
			if(IN_DATA(56) < IN_DATA(57)) begin
				TEMP_EVEN(29) = IN_DATA(56);
				IN_DATA(56) = IN_DATA(57);
				IN_DATA(57) = TEMP_EVEN(29);
			end
			else begin
				TEMP_EVEN(29) = 'd0;
			end
			if(IN_DATA(58) < IN_DATA(59)) begin
				TEMP_EVEN(30) = IN_DATA(58);
				IN_DATA(58) = IN_DATA(59);
				IN_DATA(59) = TEMP_EVEN(30);
			end
			else begin
				TEMP_EVEN(30) = 'd0;
			end
			if(IN_DATA(60) < IN_DATA(61)) begin
				TEMP_EVEN(31) = IN_DATA(60);
				IN_DATA(60) = IN_DATA(61);
				IN_DATA(61) = TEMP_EVEN(31);
			end
			else begin
				TEMP_EVEN(31) = 'd0;
			end
			if(IN_DATA(62) < IN_DATA(63)) begin
				TEMP_EVEN(32) = IN_DATA(62);
				IN_DATA(62) = IN_DATA(63);
				IN_DATA(63) = TEMP_EVEN(32);
			end
			else begin
				TEMP_EVEN(32) = 'd0;
			end
			if(IN_DATA(64) < IN_DATA(65)) begin
				TEMP_EVEN(33) = IN_DATA(64);
				IN_DATA(64) = IN_DATA(65);
				IN_DATA(65) = TEMP_EVEN(33);
			end
			else begin
				TEMP_EVEN(33) = 'd0;
			end
			if(IN_DATA(66) < IN_DATA(67)) begin
				TEMP_EVEN(34) = IN_DATA(66);
				IN_DATA(66) = IN_DATA(67);
				IN_DATA(67) = TEMP_EVEN(34);
			end
			else begin
				TEMP_EVEN(34) = 'd0;
			end
			if(IN_DATA(68) < IN_DATA(69)) begin
				TEMP_EVEN(35) = IN_DATA(68);
				IN_DATA(68) = IN_DATA(69);
				IN_DATA(69) = TEMP_EVEN(35);
			end
			else begin
				TEMP_EVEN(35) = 'd0;
			end
			if(IN_DATA(70) < IN_DATA(71)) begin
				TEMP_EVEN(36) = IN_DATA(70);
				IN_DATA(70) = IN_DATA(71);
				IN_DATA(71) = TEMP_EVEN(36);
			end
			else begin
				TEMP_EVEN(36) = 'd0;
			end
			if(IN_DATA(72) < IN_DATA(73)) begin
				TEMP_EVEN(37) = IN_DATA(72);
				IN_DATA(72) = IN_DATA(73);
				IN_DATA(73) = TEMP_EVEN(37);
			end
			else begin
				TEMP_EVEN(37) = 'd0;
			end
			if(IN_DATA(74) < IN_DATA(75)) begin
				TEMP_EVEN(38) = IN_DATA(74);
				IN_DATA(74) = IN_DATA(75);
				IN_DATA(75) = TEMP_EVEN(38);
			end
			else begin
				TEMP_EVEN(38) = 'd0;
			end
			if(IN_DATA(76) < IN_DATA(77)) begin
				TEMP_EVEN(39) = IN_DATA(76);
				IN_DATA(76) = IN_DATA(77);
				IN_DATA(77) = TEMP_EVEN(39);
			end
			else begin
				TEMP_EVEN(39) = 'd0;
			end
			if(IN_DATA(78) < IN_DATA(79)) begin
				TEMP_EVEN(40) = IN_DATA(78);
				IN_DATA(78) = IN_DATA(79);
				IN_DATA(79) = TEMP_EVEN(40);
			end
			else begin
				TEMP_EVEN(40) = 'd0;
			end
			if(IN_DATA(80) < IN_DATA(81)) begin
				TEMP_EVEN(41) = IN_DATA(80);
				IN_DATA(80) = IN_DATA(81);
				IN_DATA(81) = TEMP_EVEN(41);
			end
			else begin
				TEMP_EVEN(41) = 'd0;
			end
			if(IN_DATA(82) < IN_DATA(83)) begin
				TEMP_EVEN(42) = IN_DATA(82);
				IN_DATA(82) = IN_DATA(83);
				IN_DATA(83) = TEMP_EVEN(42);
			end
			else begin
				TEMP_EVEN(42) = 'd0;
			end
			if(IN_DATA(84) < IN_DATA(85)) begin
				TEMP_EVEN(43) = IN_DATA(84);
				IN_DATA(84) = IN_DATA(85);
				IN_DATA(85) = TEMP_EVEN(43);
			end
			else begin
				TEMP_EVEN(43) = 'd0;
			end
			if(IN_DATA(86) < IN_DATA(87)) begin
				TEMP_EVEN(44) = IN_DATA(86);
				IN_DATA(86) = IN_DATA(87);
				IN_DATA(87) = TEMP_EVEN(44);
			end
			else begin
				TEMP_EVEN(44) = 'd0;
			end
			if(IN_DATA(88) < IN_DATA(89)) begin
				TEMP_EVEN(45) = IN_DATA(88);
				IN_DATA(88) = IN_DATA(89);
				IN_DATA(89) = TEMP_EVEN(45);
			end
			else begin
				TEMP_EVEN(45) = 'd0;
			end
			if(IN_DATA(90) < IN_DATA(91)) begin
				TEMP_EVEN(46) = IN_DATA(90);
				IN_DATA(90) = IN_DATA(91);
				IN_DATA(91) = TEMP_EVEN(46);
			end
			else begin
				TEMP_EVEN(46) = 'd0;
			end
			if(IN_DATA(92) < IN_DATA(93)) begin
				TEMP_EVEN(47) = IN_DATA(92);
				IN_DATA(92) = IN_DATA(93);
				IN_DATA(93) = TEMP_EVEN(47);
			end
			else begin
				TEMP_EVEN(47) = 'd0;
			end
			if(IN_DATA(94) < IN_DATA(95)) begin
				TEMP_EVEN(48) = IN_DATA(94);
				IN_DATA(94) = IN_DATA(95);
				IN_DATA(95) = TEMP_EVEN(48);
			end
			else begin
				TEMP_EVEN(48) = 'd0;
			end
			if(IN_DATA(96) < IN_DATA(97)) begin
				TEMP_EVEN(49) = IN_DATA(96);
				IN_DATA(96) = IN_DATA(97);
				IN_DATA(97) = TEMP_EVEN(49);
			end
			else begin
				TEMP_EVEN(49) = 'd0;
			end
			if(IN_DATA(98) < IN_DATA(99)) begin
				TEMP_EVEN(50) = IN_DATA(98);
				IN_DATA(98) = IN_DATA(99);
				IN_DATA(99) = TEMP_EVEN(50);
			end
			else begin
				TEMP_EVEN(50) = 'd0;
			end
			if(IN_DATA(100) < IN_DATA(101)) begin
				TEMP_EVEN(51) = IN_DATA(100);
				IN_DATA(100) = IN_DATA(101);
				IN_DATA(101) = TEMP_EVEN(51);
			end
			else begin
				TEMP_EVEN(51) = 'd0;
			end
			if(IN_DATA(102) < IN_DATA(103)) begin
				TEMP_EVEN(52) = IN_DATA(102);
				IN_DATA(102) = IN_DATA(103);
				IN_DATA(103) = TEMP_EVEN(52);
			end
			else begin
				TEMP_EVEN(52) = 'd0;
			end
			if(IN_DATA(104) < IN_DATA(105)) begin
				TEMP_EVEN(53) = IN_DATA(104);
				IN_DATA(104) = IN_DATA(105);
				IN_DATA(105) = TEMP_EVEN(53);
			end
			else begin
				TEMP_EVEN(53) = 'd0;
			end
			if(IN_DATA(106) < IN_DATA(107)) begin
				TEMP_EVEN(54) = IN_DATA(106);
				IN_DATA(106) = IN_DATA(107);
				IN_DATA(107) = TEMP_EVEN(54);
			end
			else begin
				TEMP_EVEN(54) = 'd0;
			end
			if(IN_DATA(108) < IN_DATA(109)) begin
				TEMP_EVEN(55) = IN_DATA(108);
				IN_DATA(108) = IN_DATA(109);
				IN_DATA(109) = TEMP_EVEN(55);
			end
			else begin
				TEMP_EVEN(55) = 'd0;
			end
			if(IN_DATA(110) < IN_DATA(111)) begin
				TEMP_EVEN(56) = IN_DATA(110);
				IN_DATA(110) = IN_DATA(111);
				IN_DATA(111) = TEMP_EVEN(56);
			end
			else begin
				TEMP_EVEN(56) = 'd0;
			end
			if(IN_DATA(112) < IN_DATA(113)) begin
				TEMP_EVEN(57) = IN_DATA(112);
				IN_DATA(112) = IN_DATA(113);
				IN_DATA(113) = TEMP_EVEN(57);
			end
			else begin
				TEMP_EVEN(57) = 'd0;
			end
			if(IN_DATA(114) < IN_DATA(115)) begin
				TEMP_EVEN(58) = IN_DATA(114);
				IN_DATA(114) = IN_DATA(115);
				IN_DATA(115) = TEMP_EVEN(58);
			end
			else begin
				TEMP_EVEN(58) = 'd0;
			end
			if(IN_DATA(116) < IN_DATA(117)) begin
				TEMP_EVEN(59) = IN_DATA(116);
				IN_DATA(116) = IN_DATA(117);
				IN_DATA(117) = TEMP_EVEN(59);
			end
			else begin
				TEMP_EVEN(59) = 'd0;
			end
			if(IN_DATA(118) < IN_DATA(119)) begin
				TEMP_EVEN(60) = IN_DATA(118);
				IN_DATA(118) = IN_DATA(119);
				IN_DATA(119) = TEMP_EVEN(60);
			end
			else begin
				TEMP_EVEN(60) = 'd0;
			end
			if(IN_DATA(120) < IN_DATA(121)) begin
				TEMP_EVEN(61) = IN_DATA(120);
				IN_DATA(120) = IN_DATA(121);
				IN_DATA(121) = TEMP_EVEN(61);
			end
			else begin
				TEMP_EVEN(61) = 'd0;
			end
			if(IN_DATA(122) < IN_DATA(123)) begin
				TEMP_EVEN(62) = IN_DATA(122);
				IN_DATA(122) = IN_DATA(123);
				IN_DATA(123) = TEMP_EVEN(62);
			end
			else begin
				TEMP_EVEN(62) = 'd0;
			end
			if(IN_DATA(124) < IN_DATA(125)) begin
				TEMP_EVEN(63) = IN_DATA(124);
				IN_DATA(124) = IN_DATA(125);
				IN_DATA(125) = TEMP_EVEN(63);
			end
			else begin
				TEMP_EVEN(63) = 'd0;
			end
			if(IN_DATA(126) < IN_DATA(127)) begin
				TEMP_EVEN(64) = IN_DATA(126);
				IN_DATA(126) = IN_DATA(127);
				IN_DATA(127) = TEMP_EVEN(64);
			end
			else begin
				TEMP_EVEN(64) = 'd0;
			end
			if(IN_DATA(128) < IN_DATA(129)) begin
				TEMP_EVEN(65) = IN_DATA(128);
				IN_DATA(128) = IN_DATA(129);
				IN_DATA(129) = TEMP_EVEN(65);
			end
			else begin
				TEMP_EVEN(65) = 'd0;
			end
			if(IN_DATA(130) < IN_DATA(131)) begin
				TEMP_EVEN(66) = IN_DATA(130);
				IN_DATA(130) = IN_DATA(131);
				IN_DATA(131) = TEMP_EVEN(66);
			end
			else begin
				TEMP_EVEN(66) = 'd0;
			end
			if(IN_DATA(132) < IN_DATA(133)) begin
				TEMP_EVEN(67) = IN_DATA(132);
				IN_DATA(132) = IN_DATA(133);
				IN_DATA(133) = TEMP_EVEN(67);
			end
			else begin
				TEMP_EVEN(67) = 'd0;
			end
			if(IN_DATA(134) < IN_DATA(135)) begin
				TEMP_EVEN(68) = IN_DATA(134);
				IN_DATA(134) = IN_DATA(135);
				IN_DATA(135) = TEMP_EVEN(68);
			end
			else begin
				TEMP_EVEN(68) = 'd0;
			end
			if(IN_DATA(136) < IN_DATA(137)) begin
				TEMP_EVEN(69) = IN_DATA(136);
				IN_DATA(136) = IN_DATA(137);
				IN_DATA(137) = TEMP_EVEN(69);
			end
			else begin
				TEMP_EVEN(69) = 'd0;
			end
			if(IN_DATA(138) < IN_DATA(139)) begin
				TEMP_EVEN(70) = IN_DATA(138);
				IN_DATA(138) = IN_DATA(139);
				IN_DATA(139) = TEMP_EVEN(70);
			end
			else begin
				TEMP_EVEN(70) = 'd0;
			end
			if(IN_DATA(140) < IN_DATA(141)) begin
				TEMP_EVEN(71) = IN_DATA(140);
				IN_DATA(140) = IN_DATA(141);
				IN_DATA(141) = TEMP_EVEN(71);
			end
			else begin
				TEMP_EVEN(71) = 'd0;
			end
			if(IN_DATA(142) < IN_DATA(143)) begin
				TEMP_EVEN(72) = IN_DATA(142);
				IN_DATA(142) = IN_DATA(143);
				IN_DATA(143) = TEMP_EVEN(72);
			end
			else begin
				TEMP_EVEN(72) = 'd0;
			end
			if(IN_DATA(144) < IN_DATA(145)) begin
				TEMP_EVEN(73) = IN_DATA(144);
				IN_DATA(144) = IN_DATA(145);
				IN_DATA(145) = TEMP_EVEN(73);
			end
			else begin
				TEMP_EVEN(73) = 'd0;
			end
			if(IN_DATA(146) < IN_DATA(147)) begin
				TEMP_EVEN(74) = IN_DATA(146);
				IN_DATA(146) = IN_DATA(147);
				IN_DATA(147) = TEMP_EVEN(74);
			end
			else begin
				TEMP_EVEN(74) = 'd0;
			end
			if(IN_DATA(148) < IN_DATA(149)) begin
				TEMP_EVEN(75) = IN_DATA(148);
				IN_DATA(148) = IN_DATA(149);
				IN_DATA(149) = TEMP_EVEN(75);
			end
			else begin
				TEMP_EVEN(75) = 'd0;
			end
			if(IN_DATA(150) < IN_DATA(151)) begin
				TEMP_EVEN(76) = IN_DATA(150);
				IN_DATA(150) = IN_DATA(151);
				IN_DATA(151) = TEMP_EVEN(76);
			end
			else begin
				TEMP_EVEN(76) = 'd0;
			end
			if(IN_DATA(152) < IN_DATA(153)) begin
				TEMP_EVEN(77) = IN_DATA(152);
				IN_DATA(152) = IN_DATA(153);
				IN_DATA(153) = TEMP_EVEN(77);
			end
			else begin
				TEMP_EVEN(77) = 'd0;
			end
			if(IN_DATA(154) < IN_DATA(155)) begin
				TEMP_EVEN(78) = IN_DATA(154);
				IN_DATA(154) = IN_DATA(155);
				IN_DATA(155) = TEMP_EVEN(78);
			end
			else begin
				TEMP_EVEN(78) = 'd0;
			end
			if(IN_DATA(156) < IN_DATA(157)) begin
				TEMP_EVEN(79) = IN_DATA(156);
				IN_DATA(156) = IN_DATA(157);
				IN_DATA(157) = TEMP_EVEN(79);
			end
			else begin
				TEMP_EVEN(79) = 'd0;
			end
			if(IN_DATA(158) < IN_DATA(159)) begin
				TEMP_EVEN(80) = IN_DATA(158);
				IN_DATA(158) = IN_DATA(159);
				IN_DATA(159) = TEMP_EVEN(80);
			end
			else begin
				TEMP_EVEN(80) = 'd0;
			end
			if(IN_DATA(160) < IN_DATA(161)) begin
				TEMP_EVEN(81) = IN_DATA(160);
				IN_DATA(160) = IN_DATA(161);
				IN_DATA(161) = TEMP_EVEN(81);
			end
			else begin
				TEMP_EVEN(81) = 'd0;
			end
			if(IN_DATA(162) < IN_DATA(163)) begin
				TEMP_EVEN(82) = IN_DATA(162);
				IN_DATA(162) = IN_DATA(163);
				IN_DATA(163) = TEMP_EVEN(82);
			end
			else begin
				TEMP_EVEN(82) = 'd0;
			end
			if(IN_DATA(164) < IN_DATA(165)) begin
				TEMP_EVEN(83) = IN_DATA(164);
				IN_DATA(164) = IN_DATA(165);
				IN_DATA(165) = TEMP_EVEN(83);
			end
			else begin
				TEMP_EVEN(83) = 'd0;
			end
			if(IN_DATA(166) < IN_DATA(167)) begin
				TEMP_EVEN(84) = IN_DATA(166);
				IN_DATA(166) = IN_DATA(167);
				IN_DATA(167) = TEMP_EVEN(84);
			end
			else begin
				TEMP_EVEN(84) = 'd0;
			end
			if(IN_DATA(168) < IN_DATA(169)) begin
				TEMP_EVEN(85) = IN_DATA(168);
				IN_DATA(168) = IN_DATA(169);
				IN_DATA(169) = TEMP_EVEN(85);
			end
			else begin
				TEMP_EVEN(85) = 'd0;
			end
			if(IN_DATA(170) < IN_DATA(171)) begin
				TEMP_EVEN(86) = IN_DATA(170);
				IN_DATA(170) = IN_DATA(171);
				IN_DATA(171) = TEMP_EVEN(86);
			end
			else begin
				TEMP_EVEN(86) = 'd0;
			end
			if(IN_DATA(172) < IN_DATA(173)) begin
				TEMP_EVEN(87) = IN_DATA(172);
				IN_DATA(172) = IN_DATA(173);
				IN_DATA(173) = TEMP_EVEN(87);
			end
			else begin
				TEMP_EVEN(87) = 'd0;
			end
			if(IN_DATA(174) < IN_DATA(175)) begin
				TEMP_EVEN(88) = IN_DATA(174);
				IN_DATA(174) = IN_DATA(175);
				IN_DATA(175) = TEMP_EVEN(88);
			end
			else begin
				TEMP_EVEN(88) = 'd0;
			end
			if(IN_DATA(176) < IN_DATA(177)) begin
				TEMP_EVEN(89) = IN_DATA(176);
				IN_DATA(176) = IN_DATA(177);
				IN_DATA(177) = TEMP_EVEN(89);
			end
			else begin
				TEMP_EVEN(89) = 'd0;
			end
			if(IN_DATA(178) < IN_DATA(179)) begin
				TEMP_EVEN(90) = IN_DATA(178);
				IN_DATA(178) = IN_DATA(179);
				IN_DATA(179) = TEMP_EVEN(90);
			end
			else begin
				TEMP_EVEN(90) = 'd0;
			end
			if(IN_DATA(180) < IN_DATA(181)) begin
				TEMP_EVEN(91) = IN_DATA(180);
				IN_DATA(180) = IN_DATA(181);
				IN_DATA(181) = TEMP_EVEN(91);
			end
			else begin
				TEMP_EVEN(91) = 'd0;
			end
			if(IN_DATA(182) < IN_DATA(183)) begin
				TEMP_EVEN(92) = IN_DATA(182);
				IN_DATA(182) = IN_DATA(183);
				IN_DATA(183) = TEMP_EVEN(92);
			end
			else begin
				TEMP_EVEN(92) = 'd0;
			end
			if(IN_DATA(184) < IN_DATA(185)) begin
				TEMP_EVEN(93) = IN_DATA(184);
				IN_DATA(184) = IN_DATA(185);
				IN_DATA(185) = TEMP_EVEN(93);
			end
			else begin
				TEMP_EVEN(93) = 'd0;
			end
			if(IN_DATA(186) < IN_DATA(187)) begin
				TEMP_EVEN(94) = IN_DATA(186);
				IN_DATA(186) = IN_DATA(187);
				IN_DATA(187) = TEMP_EVEN(94);
			end
			else begin
				TEMP_EVEN(94) = 'd0;
			end
			if(IN_DATA(188) < IN_DATA(189)) begin
				TEMP_EVEN(95) = IN_DATA(188);
				IN_DATA(188) = IN_DATA(189);
				IN_DATA(189) = TEMP_EVEN(95);
			end
			else begin
				TEMP_EVEN(95) = 'd0;
			end
			if(IN_DATA(190) < IN_DATA(191)) begin
				TEMP_EVEN(96) = IN_DATA(190);
				IN_DATA(190) = IN_DATA(191);
				IN_DATA(191) = TEMP_EVEN(96);
			end
			else begin
				TEMP_EVEN(96) = 'd0;
			end
			if(IN_DATA(192) < IN_DATA(193)) begin
				TEMP_EVEN(97) = IN_DATA(192);
				IN_DATA(192) = IN_DATA(193);
				IN_DATA(193) = TEMP_EVEN(97);
			end
			else begin
				TEMP_EVEN(97) = 'd0;
			end
			if(IN_DATA(194) < IN_DATA(195)) begin
				TEMP_EVEN(98) = IN_DATA(194);
				IN_DATA(194) = IN_DATA(195);
				IN_DATA(195) = TEMP_EVEN(98);
			end
			else begin
				TEMP_EVEN(98) = 'd0;
			end
			if(IN_DATA(196) < IN_DATA(197)) begin
				TEMP_EVEN(99) = IN_DATA(196);
				IN_DATA(196) = IN_DATA(197);
				IN_DATA(197) = TEMP_EVEN(99);
			end
			else begin
				TEMP_EVEN(99) = 'd0;
			end
			if(IN_DATA(198) < IN_DATA(199)) begin
				TEMP_EVEN(100) = IN_DATA(198);
				IN_DATA(198) = IN_DATA(199);
				IN_DATA(199) = TEMP_EVEN(100);
			end
			else begin
				TEMP_EVEN(100) = 'd0;
			end
			if(IN_DATA(200) < IN_DATA(201)) begin
				TEMP_EVEN(101) = IN_DATA(200);
				IN_DATA(200) = IN_DATA(201);
				IN_DATA(201) = TEMP_EVEN(101);
			end
			else begin
				TEMP_EVEN(101) = 'd0;
			end
			if(IN_DATA(202) < IN_DATA(203)) begin
				TEMP_EVEN(102) = IN_DATA(202);
				IN_DATA(202) = IN_DATA(203);
				IN_DATA(203) = TEMP_EVEN(102);
			end
			else begin
				TEMP_EVEN(102) = 'd0;
			end
			if(IN_DATA(204) < IN_DATA(205)) begin
				TEMP_EVEN(103) = IN_DATA(204);
				IN_DATA(204) = IN_DATA(205);
				IN_DATA(205) = TEMP_EVEN(103);
			end
			else begin
				TEMP_EVEN(103) = 'd0;
			end
			if(IN_DATA(206) < IN_DATA(207)) begin
				TEMP_EVEN(104) = IN_DATA(206);
				IN_DATA(206) = IN_DATA(207);
				IN_DATA(207) = TEMP_EVEN(104);
			end
			else begin
				TEMP_EVEN(104) = 'd0;
			end
			if(IN_DATA(208) < IN_DATA(209)) begin
				TEMP_EVEN(105) = IN_DATA(208);
				IN_DATA(208) = IN_DATA(209);
				IN_DATA(209) = TEMP_EVEN(105);
			end
			else begin
				TEMP_EVEN(105) = 'd0;
			end
			if(IN_DATA(210) < IN_DATA(211)) begin
				TEMP_EVEN(106) = IN_DATA(210);
				IN_DATA(210) = IN_DATA(211);
				IN_DATA(211) = TEMP_EVEN(106);
			end
			else begin
				TEMP_EVEN(106) = 'd0;
			end
			if(IN_DATA(212) < IN_DATA(213)) begin
				TEMP_EVEN(107) = IN_DATA(212);
				IN_DATA(212) = IN_DATA(213);
				IN_DATA(213) = TEMP_EVEN(107);
			end
			else begin
				TEMP_EVEN(107) = 'd0;
			end
			if(IN_DATA(214) < IN_DATA(215)) begin
				TEMP_EVEN(108) = IN_DATA(214);
				IN_DATA(214) = IN_DATA(215);
				IN_DATA(215) = TEMP_EVEN(108);
			end
			else begin
				TEMP_EVEN(108) = 'd0;
			end
			if(IN_DATA(216) < IN_DATA(217)) begin
				TEMP_EVEN(109) = IN_DATA(216);
				IN_DATA(216) = IN_DATA(217);
				IN_DATA(217) = TEMP_EVEN(109);
			end
			else begin
				TEMP_EVEN(109) = 'd0;
			end
			if(IN_DATA(218) < IN_DATA(219)) begin
				TEMP_EVEN(110) = IN_DATA(218);
				IN_DATA(218) = IN_DATA(219);
				IN_DATA(219) = TEMP_EVEN(110);
			end
			else begin
				TEMP_EVEN(110) = 'd0;
			end
			if(IN_DATA(220) < IN_DATA(221)) begin
				TEMP_EVEN(111) = IN_DATA(220);
				IN_DATA(220) = IN_DATA(221);
				IN_DATA(221) = TEMP_EVEN(111);
			end
			else begin
				TEMP_EVEN(111) = 'd0;
			end
			if(IN_DATA(222) < IN_DATA(223)) begin
				TEMP_EVEN(112) = IN_DATA(222);
				IN_DATA(222) = IN_DATA(223);
				IN_DATA(223) = TEMP_EVEN(112);
			end
			else begin
				TEMP_EVEN(112) = 'd0;
			end
			if(IN_DATA(224) < IN_DATA(225)) begin
				TEMP_EVEN(113) = IN_DATA(224);
				IN_DATA(224) = IN_DATA(225);
				IN_DATA(225) = TEMP_EVEN(113);
			end
			else begin
				TEMP_EVEN(113) = 'd0;
			end
			if(IN_DATA(226) < IN_DATA(227)) begin
				TEMP_EVEN(114) = IN_DATA(226);
				IN_DATA(226) = IN_DATA(227);
				IN_DATA(227) = TEMP_EVEN(114);
			end
			else begin
				TEMP_EVEN(114) = 'd0;
			end
			if(IN_DATA(228) < IN_DATA(229)) begin
				TEMP_EVEN(115) = IN_DATA(228);
				IN_DATA(228) = IN_DATA(229);
				IN_DATA(229) = TEMP_EVEN(115);
			end
			else begin
				TEMP_EVEN(115) = 'd0;
			end
			if(IN_DATA(230) < IN_DATA(231)) begin
				TEMP_EVEN(116) = IN_DATA(230);
				IN_DATA(230) = IN_DATA(231);
				IN_DATA(231) = TEMP_EVEN(116);
			end
			else begin
				TEMP_EVEN(116) = 'd0;
			end
			if(IN_DATA(232) < IN_DATA(233)) begin
				TEMP_EVEN(117) = IN_DATA(232);
				IN_DATA(232) = IN_DATA(233);
				IN_DATA(233) = TEMP_EVEN(117);
			end
			else begin
				TEMP_EVEN(117) = 'd0;
			end
			if(IN_DATA(234) < IN_DATA(235)) begin
				TEMP_EVEN(118) = IN_DATA(234);
				IN_DATA(234) = IN_DATA(235);
				IN_DATA(235) = TEMP_EVEN(118);
			end
			else begin
				TEMP_EVEN(118) = 'd0;
			end
			if(IN_DATA(236) < IN_DATA(237)) begin
				TEMP_EVEN(119) = IN_DATA(236);
				IN_DATA(236) = IN_DATA(237);
				IN_DATA(237) = TEMP_EVEN(119);
			end
			else begin
				TEMP_EVEN(119) = 'd0;
			end
			if(IN_DATA(238) < IN_DATA(239)) begin
				TEMP_EVEN(120) = IN_DATA(238);
				IN_DATA(238) = IN_DATA(239);
				IN_DATA(239) = TEMP_EVEN(120);
			end
			else begin
				TEMP_EVEN(120) = 'd0;
			end
			if(IN_DATA(240) < IN_DATA(241)) begin
				TEMP_EVEN(121) = IN_DATA(240);
				IN_DATA(240) = IN_DATA(241);
				IN_DATA(241) = TEMP_EVEN(121);
			end
			else begin
				TEMP_EVEN(121) = 'd0;
			end
			if(IN_DATA(242) < IN_DATA(243)) begin
				TEMP_EVEN(122) = IN_DATA(242);
				IN_DATA(242) = IN_DATA(243);
				IN_DATA(243) = TEMP_EVEN(122);
			end
			else begin
				TEMP_EVEN(122) = 'd0;
			end
			if(IN_DATA(244) < IN_DATA(245)) begin
				TEMP_EVEN(123) = IN_DATA(244);
				IN_DATA(244) = IN_DATA(245);
				IN_DATA(245) = TEMP_EVEN(123);
			end
			else begin
				TEMP_EVEN(123) = 'd0;
			end
			if(IN_DATA(246) < IN_DATA(247)) begin
				TEMP_EVEN(124) = IN_DATA(246);
				IN_DATA(246) = IN_DATA(247);
				IN_DATA(247) = TEMP_EVEN(124);
			end
			else begin
				TEMP_EVEN(124) = 'd0;
			end
			if(IN_DATA(248) < IN_DATA(249)) begin
				TEMP_EVEN(125) = IN_DATA(248);
				IN_DATA(248) = IN_DATA(249);
				IN_DATA(249) = TEMP_EVEN(125);
			end
			else begin
				TEMP_EVEN(125) = 'd0;
			end
			if(IN_DATA(250) < IN_DATA(251)) begin
				TEMP_EVEN(126) = IN_DATA(250);
				IN_DATA(250) = IN_DATA(251);
				IN_DATA(251) = TEMP_EVEN(126);
			end
			else begin
				TEMP_EVEN(126) = 'd0;
			end
			if(IN_DATA(252) < IN_DATA(253)) begin
				TEMP_EVEN(127) = IN_DATA(252);
				IN_DATA(252) = IN_DATA(253);
				IN_DATA(253) = TEMP_EVEN(127);
			end
			else begin
				TEMP_EVEN(127) = 'd0;
			end
			if(IN_DATA(254) < IN_DATA(255)) begin
				TEMP_EVEN(128) = IN_DATA(254);
				IN_DATA(254) = IN_DATA(255);
				IN_DATA(255) = TEMP_EVEN(128);
			end
			else begin
				TEMP_EVEN(128) = 'd0;
			end
		end
	end
	else begin
		TEMP_ODD(0) = 'd0;
		TEMP_ODD(1) = 'd0;
		TEMP_ODD(2) = 'd0;
		TEMP_ODD(3) = 'd0;
		TEMP_ODD(4) = 'd0;
		TEMP_ODD(5) = 'd0;
		TEMP_ODD(6) = 'd0;
		TEMP_ODD(7) = 'd0;
		TEMP_ODD(8) = 'd0;
		TEMP_ODD(9) = 'd0;
		TEMP_ODD(10) = 'd0;
		TEMP_ODD(11) = 'd0;
		TEMP_ODD(12) = 'd0;
		TEMP_ODD(13) = 'd0;
		TEMP_ODD(14) = 'd0;
		TEMP_ODD(15) = 'd0;
		TEMP_ODD(16) = 'd0;
		TEMP_ODD(17) = 'd0;
		TEMP_ODD(18) = 'd0;
		TEMP_ODD(19) = 'd0;
		TEMP_ODD(20) = 'd0;
		TEMP_ODD(21) = 'd0;
		TEMP_ODD(22) = 'd0;
		TEMP_ODD(23) = 'd0;
		TEMP_ODD(24) = 'd0;
		TEMP_ODD(25) = 'd0;
		TEMP_ODD(26) = 'd0;
		TEMP_ODD(27) = 'd0;
		TEMP_ODD(28) = 'd0;
		TEMP_ODD(29) = 'd0;
		TEMP_ODD(30) = 'd0;
		TEMP_ODD(31) = 'd0;
		TEMP_ODD(32) = 'd0;
		TEMP_ODD(33) = 'd0;
		TEMP_ODD(34) = 'd0;
		TEMP_ODD(35) = 'd0;
		TEMP_ODD(36) = 'd0;
		TEMP_ODD(37) = 'd0;
		TEMP_ODD(38) = 'd0;
		TEMP_ODD(39) = 'd0;
		TEMP_ODD(40) = 'd0;
		TEMP_ODD(41) = 'd0;
		TEMP_ODD(42) = 'd0;
		TEMP_ODD(43) = 'd0;
		TEMP_ODD(44) = 'd0;
		TEMP_ODD(45) = 'd0;
		TEMP_ODD(46) = 'd0;
		TEMP_ODD(47) = 'd0;
		TEMP_ODD(48) = 'd0;
		TEMP_ODD(49) = 'd0;
		TEMP_ODD(50) = 'd0;
		TEMP_ODD(51) = 'd0;
		TEMP_ODD(52) = 'd0;
		TEMP_ODD(53) = 'd0;
		TEMP_ODD(54) = 'd0;
		TEMP_ODD(55) = 'd0;
		TEMP_ODD(56) = 'd0;
		TEMP_ODD(57) = 'd0;
		TEMP_ODD(58) = 'd0;
		TEMP_ODD(59) = 'd0;
		TEMP_ODD(60) = 'd0;
		TEMP_ODD(61) = 'd0;
		TEMP_ODD(62) = 'd0;
		TEMP_ODD(63) = 'd0;
		TEMP_ODD(64) = 'd0;
		TEMP_ODD(65) = 'd0;
		TEMP_ODD(66) = 'd0;
		TEMP_ODD(67) = 'd0;
		TEMP_ODD(68) = 'd0;
		TEMP_ODD(69) = 'd0;
		TEMP_ODD(70) = 'd0;
		TEMP_ODD(71) = 'd0;
		TEMP_ODD(72) = 'd0;
		TEMP_ODD(73) = 'd0;
		TEMP_ODD(74) = 'd0;
		TEMP_ODD(75) = 'd0;
		TEMP_ODD(76) = 'd0;
		TEMP_ODD(77) = 'd0;
		TEMP_ODD(78) = 'd0;
		TEMP_ODD(79) = 'd0;
		TEMP_ODD(80) = 'd0;
		TEMP_ODD(81) = 'd0;
		TEMP_ODD(82) = 'd0;
		TEMP_ODD(83) = 'd0;
		TEMP_ODD(84) = 'd0;
		TEMP_ODD(85) = 'd0;
		TEMP_ODD(86) = 'd0;
		TEMP_ODD(87) = 'd0;
		TEMP_ODD(88) = 'd0;
		TEMP_ODD(89) = 'd0;
		TEMP_ODD(90) = 'd0;
		TEMP_ODD(91) = 'd0;
		TEMP_ODD(92) = 'd0;
		TEMP_ODD(93) = 'd0;
		TEMP_ODD(94) = 'd0;
		TEMP_ODD(95) = 'd0;
		TEMP_ODD(96) = 'd0;
		TEMP_ODD(97) = 'd0;
		TEMP_ODD(98) = 'd0;
		TEMP_ODD(99) = 'd0;
		TEMP_ODD(100) = 'd0;
		TEMP_ODD(101) = 'd0;
		TEMP_ODD(102) = 'd0;
		TEMP_ODD(103) = 'd0;
		TEMP_ODD(104) = 'd0;
		TEMP_ODD(105) = 'd0;
		TEMP_ODD(106) = 'd0;
		TEMP_ODD(107) = 'd0;
		TEMP_ODD(108) = 'd0;
		TEMP_ODD(109) = 'd0;
		TEMP_ODD(110) = 'd0;
		TEMP_ODD(111) = 'd0;
		TEMP_ODD(112) = 'd0;
		TEMP_ODD(113) = 'd0;
		TEMP_ODD(114) = 'd0;
		TEMP_ODD(115) = 'd0;
		TEMP_ODD(116) = 'd0;
		TEMP_ODD(117) = 'd0;
		TEMP_ODD(118) = 'd0;
		TEMP_ODD(119) = 'd0;
		TEMP_ODD(120) = 'd0;
		TEMP_ODD(120) = 'd0;
		TEMP_ODD(121) = 'd0;
		TEMP_ODD(122) = 'd0;
		TEMP_ODD(123) = 'd0;
		TEMP_ODD(124) = 'd0;
		TEMP_ODD(125) = 'd0;
		TEMP_ODD(126) = 'd0;
		TEMP_ODD(127) = 'd0;

		TEMP_EVEN(0) = 'd0;
		TEMP_EVEN(1) = 'd0;
		TEMP_EVEN(2) = 'd0;
		TEMP_EVEN(3) = 'd0;
		TEMP_EVEN(4) = 'd0;
		TEMP_EVEN(5) = 'd0;
		TEMP_EVEN(6) = 'd0;
		TEMP_EVEN(7) = 'd0;
		TEMP_EVEN(8) = 'd0;
		TEMP_EVEN(9) = 'd0;
		TEMP_EVEN(10) = 'd0;
		TEMP_EVEN(11) = 'd0;
		TEMP_EVEN(12) = 'd0;
		TEMP_EVEN(13) = 'd0;
		TEMP_EVEN(14) = 'd0;
		TEMP_EVEN(15) = 'd0;
		TEMP_EVEN(16) = 'd0;
		TEMP_EVEN(17) = 'd0;
		TEMP_EVEN(18) = 'd0;
		TEMP_EVEN(19) = 'd0;
		TEMP_EVEN(20) = 'd0;
		TEMP_EVEN(21) = 'd0;
		TEMP_EVEN(22) = 'd0;
		TEMP_EVEN(23) = 'd0;
		TEMP_EVEN(24) = 'd0;
		TEMP_EVEN(25) = 'd0;
		TEMP_EVEN(26) = 'd0;
		TEMP_EVEN(27) = 'd0;
		TEMP_EVEN(28) = 'd0;
		TEMP_EVEN(29) = 'd0;
		TEMP_EVEN(30) = 'd0;
		TEMP_EVEN(31) = 'd0;
		TEMP_EVEN(32) = 'd0;
		TEMP_EVEN(33) = 'd0;
		TEMP_EVEN(34) = 'd0;
		TEMP_EVEN(35) = 'd0;
		TEMP_EVEN(36) = 'd0;
		TEMP_EVEN(37) = 'd0;
		TEMP_EVEN(38) = 'd0;
		TEMP_EVEN(39) = 'd0;
		TEMP_EVEN(40) = 'd0;
		TEMP_EVEN(41) = 'd0;
		TEMP_EVEN(42) = 'd0;
		TEMP_EVEN(43) = 'd0;
		TEMP_EVEN(44) = 'd0;
		TEMP_EVEN(45) = 'd0;
		TEMP_EVEN(46) = 'd0;
		TEMP_EVEN(47) = 'd0;
		TEMP_EVEN(48) = 'd0;
		TEMP_EVEN(49) = 'd0;
		TEMP_EVEN(50) = 'd0;
		TEMP_EVEN(51) = 'd0;
		TEMP_EVEN(52) = 'd0;
		TEMP_EVEN(53) = 'd0;
		TEMP_EVEN(54) = 'd0;
		TEMP_EVEN(55) = 'd0;
		TEMP_EVEN(56) = 'd0;
		TEMP_EVEN(57) = 'd0;
		TEMP_EVEN(58) = 'd0;
		TEMP_EVEN(59) = 'd0;
		TEMP_EVEN(60) = 'd0;
		TEMP_EVEN(61) = 'd0;
		TEMP_EVEN(62) = 'd0;
		TEMP_EVEN(63) = 'd0;
		TEMP_EVEN(64) = 'd0;
		TEMP_EVEN(65) = 'd0;
		TEMP_EVEN(66) = 'd0;
		TEMP_EVEN(67) = 'd0;
		TEMP_EVEN(68) = 'd0;
		TEMP_EVEN(69) = 'd0;
		TEMP_EVEN(70) = 'd0;
		TEMP_EVEN(71) = 'd0;
		TEMP_EVEN(72) = 'd0;
		TEMP_EVEN(73) = 'd0;
		TEMP_EVEN(74) = 'd0;
		TEMP_EVEN(75) = 'd0;
		TEMP_EVEN(76) = 'd0;
		TEMP_EVEN(77) = 'd0;
		TEMP_EVEN(78) = 'd0;
		TEMP_EVEN(79) = 'd0;
		TEMP_EVEN(80) = 'd0;
		TEMP_EVEN(81) = 'd0;
		TEMP_EVEN(82) = 'd0;
		TEMP_EVEN(83) = 'd0;
		TEMP_EVEN(84) = 'd0;
		TEMP_EVEN(85) = 'd0;
		TEMP_EVEN(86) = 'd0;
		TEMP_EVEN(87) = 'd0;
		TEMP_EVEN(88) = 'd0;
		TEMP_EVEN(89) = 'd0;
		TEMP_EVEN(90) = 'd0;
		TEMP_EVEN(91) = 'd0;
		TEMP_EVEN(92) = 'd0;
		TEMP_EVEN(93) = 'd0;
		TEMP_EVEN(94) = 'd0;
		TEMP_EVEN(95) = 'd0;
		TEMP_EVEN(96) = 'd0;
		TEMP_EVEN(97) = 'd0;
		TEMP_EVEN(98) = 'd0;
		TEMP_EVEN(99) = 'd0;
		TEMP_EVEN(100) = 'd0;
		TEMP_EVEN(101) = 'd0;
		TEMP_EVEN(102) = 'd0;
		TEMP_EVEN(103) = 'd0;
		TEMP_EVEN(104) = 'd0;
		TEMP_EVEN(105) = 'd0;
		TEMP_EVEN(106) = 'd0;
		TEMP_EVEN(107) = 'd0;
		TEMP_EVEN(108) = 'd0;
		TEMP_EVEN(109) = 'd0;
		TEMP_EVEN(110) = 'd0;
		TEMP_EVEN(111) = 'd0;
		TEMP_EVEN(112) = 'd0;
		TEMP_EVEN(113) = 'd0;
		TEMP_EVEN(114) = 'd0;
		TEMP_EVEN(115) = 'd0;
		TEMP_EVEN(116) = 'd0;
		TEMP_EVEN(117) = 'd0;
		TEMP_EVEN(118) = 'd0;
		TEMP_EVEN(119) = 'd0;
		TEMP_EVEN(120) = 'd0;
		TEMP_EVEN(120) = 'd0;
		TEMP_EVEN(121) = 'd0;
		TEMP_EVEN(122) = 'd0;
		TEMP_EVEN(123) = 'd0;
		TEMP_EVEN(124) = 'd0;
		TEMP_EVEN(125) = 'd0;
		TEMP_EVEN(126) = 'd0;
		TEMP_EVEN(127) = 'd0;
		TEMP_EVEN(128) = 'd0;
	end
end

endmodule