`timescale 1ns/10ps

module Bubble_Sort(
	clk,
	rst_n,
	in_valid,
	in_data,
	out_valid,
	out_data
	);

input             clk;
input             rst_n;
input             in_valid;
input       [7:0] in_data;
output reg	      out_valid;
output reg	[7:0] out_data;

reg				  dump_out_flag;



/*
 * Memory to store in data
 */
reg			[7:0] in_data0;
reg			[7:0] in_data1;
reg			[7:0] in_data2;
reg			[7:0] in_data3;
reg			[7:0] in_data4;
reg			[7:0] in_data5;
reg			[7:0] in_data6;
reg			[7:0] in_data7;
reg			[7:0] in_data8;
reg			[7:0] in_data9;
reg			[7:0] in_data10;
reg			[7:0] in_data11;
reg			[7:0] in_data12;
reg			[7:0] in_data13;
reg			[7:0] in_data14;
reg			[7:0] in_data15;
reg			[7:0] in_data16;
reg			[7:0] in_data17;
reg			[7:0] in_data18;
reg			[7:0] in_data19;
reg			[7:0] in_data20;
reg			[7:0] in_data21;
reg			[7:0] in_data22;
reg			[7:0] in_data23;
reg			[7:0] in_data24;
reg			[7:0] in_data25;
reg			[7:0] in_data26;
reg			[7:0] in_data27;
reg			[7:0] in_data28;
reg			[7:0] in_data29;
reg			[7:0] in_data30;
reg			[7:0] in_data31;
reg			[7:0] in_data32;
reg			[7:0] in_data33;
reg			[7:0] in_data34;
reg			[7:0] in_data35;
reg			[7:0] in_data36;
reg			[7:0] in_data37;
reg			[7:0] in_data38;
reg			[7:0] in_data39;
reg			[7:0] in_data40;
reg			[7:0] in_data41;
reg			[7:0] in_data42;
reg			[7:0] in_data43;
reg			[7:0] in_data44;
reg			[7:0] in_data45;
reg			[7:0] in_data46;
reg			[7:0] in_data47;
reg			[7:0] in_data48;
reg			[7:0] in_data49;
reg			[7:0] in_data50;
reg			[7:0] in_data51;
reg			[7:0] in_data52;
reg			[7:0] in_data53;
reg			[7:0] in_data54;
reg			[7:0] in_data55;
reg			[7:0] in_data56;
reg			[7:0] in_data57;
reg			[7:0] in_data58;
reg			[7:0] in_data59;
reg			[7:0] in_data60;
reg			[7:0] in_data61;
reg			[7:0] in_data62;
reg			[7:0] in_data63;
reg			[7:0] in_data64;
reg			[7:0] in_data65;
reg			[7:0] in_data66;
reg			[7:0] in_data67;
reg			[7:0] in_data68;
reg			[7:0] in_data69;
reg			[7:0] in_data70;
reg			[7:0] in_data71;
reg			[7:0] in_data72;
reg			[7:0] in_data73;
reg			[7:0] in_data74;
reg			[7:0] in_data75;
reg			[7:0] in_data76;
reg			[7:0] in_data77;
reg			[7:0] in_data78;
reg			[7:0] in_data79;
reg			[7:0] in_data80;
reg			[7:0] in_data81;
reg			[7:0] in_data82;
reg			[7:0] in_data83;
reg			[7:0] in_data84;
reg			[7:0] in_data85;
reg			[7:0] in_data86;
reg			[7:0] in_data87;
reg			[7:0] in_data88;
reg			[7:0] in_data89;
reg			[7:0] in_data90;
reg			[7:0] in_data91;
reg			[7:0] in_data92;
reg			[7:0] in_data93;
reg			[7:0] in_data94;
reg			[7:0] in_data95;
reg			[7:0] in_data96;
reg			[7:0] in_data97;
reg			[7:0] in_data98;
reg			[7:0] in_data99;
reg			[7:0] in_data100;
reg			[7:0] in_data101;
reg			[7:0] in_data102;
reg			[7:0] in_data103;
reg			[7:0] in_data104;
reg			[7:0] in_data105;
reg			[7:0] in_data106;
reg			[7:0] in_data107;
reg			[7:0] in_data108;
reg			[7:0] in_data109;
reg			[7:0] in_data110;
reg			[7:0] in_data111;
reg			[7:0] in_data112;
reg			[7:0] in_data113;
reg			[7:0] in_data114;
reg			[7:0] in_data115;
reg			[7:0] in_data116;
reg			[7:0] in_data117;
reg			[7:0] in_data118;
reg			[7:0] in_data119;
reg			[7:0] in_data120;
reg			[7:0] in_data121;
reg			[7:0] in_data122;
reg			[7:0] in_data123;
reg			[7:0] in_data124;
reg			[7:0] in_data125;
reg			[7:0] in_data126;
reg			[7:0] in_data127;
reg			[7:0] in_data128;
reg			[7:0] in_data129;
reg			[7:0] in_data130;
reg			[7:0] in_data131;
reg			[7:0] in_data132;
reg			[7:0] in_data133;
reg			[7:0] in_data134;
reg			[7:0] in_data135;
reg			[7:0] in_data136;
reg			[7:0] in_data137;
reg			[7:0] in_data138;
reg			[7:0] in_data139;
reg			[7:0] in_data140;
reg			[7:0] in_data141;
reg			[7:0] in_data142;
reg			[7:0] in_data143;
reg			[7:0] in_data144;
reg			[7:0] in_data145;
reg			[7:0] in_data146;
reg			[7:0] in_data147;
reg			[7:0] in_data148;
reg			[7:0] in_data149;
reg			[7:0] in_data150;
reg			[7:0] in_data151;
reg			[7:0] in_data152;
reg			[7:0] in_data153;
reg			[7:0] in_data154;
reg			[7:0] in_data155;
reg			[7:0] in_data156;
reg			[7:0] in_data157;
reg			[7:0] in_data158;
reg			[7:0] in_data159;
reg			[7:0] in_data160;
reg			[7:0] in_data161;
reg			[7:0] in_data162;
reg			[7:0] in_data163;
reg			[7:0] in_data164;
reg			[7:0] in_data165;
reg			[7:0] in_data166;
reg			[7:0] in_data167;
reg			[7:0] in_data168;
reg			[7:0] in_data169;
reg			[7:0] in_data170;
reg			[7:0] in_data171;
reg			[7:0] in_data172;
reg			[7:0] in_data173;
reg			[7:0] in_data174;
reg			[7:0] in_data175;
reg			[7:0] in_data176;
reg			[7:0] in_data177;
reg			[7:0] in_data178;
reg			[7:0] in_data179;
reg			[7:0] in_data180;
reg			[7:0] in_data181;
reg			[7:0] in_data182;
reg			[7:0] in_data183;
reg			[7:0] in_data184;
reg			[7:0] in_data185;
reg			[7:0] in_data186;
reg			[7:0] in_data187;
reg			[7:0] in_data188;
reg			[7:0] in_data189;
reg			[7:0] in_data190;
reg			[7:0] in_data191;
reg			[7:0] in_data192;
reg			[7:0] in_data193;
reg			[7:0] in_data194;
reg			[7:0] in_data195;
reg			[7:0] in_data196;
reg			[7:0] in_data197;
reg			[7:0] in_data198;
reg			[7:0] in_data199;
reg			[7:0] in_data200;
reg			[7:0] in_data201;
reg			[7:0] in_data202;
reg			[7:0] in_data203;
reg			[7:0] in_data204;
reg			[7:0] in_data205;
reg			[7:0] in_data206;
reg			[7:0] in_data207;
reg			[7:0] in_data208;
reg			[7:0] in_data209;
reg			[7:0] in_data210;
reg			[7:0] in_data211;
reg			[7:0] in_data212;
reg			[7:0] in_data213;
reg			[7:0] in_data214;
reg			[7:0] in_data215;
reg			[7:0] in_data216;
reg			[7:0] in_data217;
reg			[7:0] in_data218;
reg			[7:0] in_data219;
reg			[7:0] in_data220;
reg			[7:0] in_data221;
reg			[7:0] in_data222;
reg			[7:0] in_data223;
reg			[7:0] in_data224;
reg			[7:0] in_data225;
reg			[7:0] in_data226;
reg			[7:0] in_data227;
reg			[7:0] in_data228;
reg			[7:0] in_data229;
reg			[7:0] in_data230;
reg			[7:0] in_data231;
reg			[7:0] in_data232;
reg			[7:0] in_data233;
reg			[7:0] in_data234;
reg			[7:0] in_data235;
reg			[7:0] in_data236;
reg			[7:0] in_data237;
reg			[7:0] in_data238;
reg			[7:0] in_data239;
reg			[7:0] in_data240;
reg			[7:0] in_data241;
reg			[7:0] in_data242;
reg			[7:0] in_data243;
reg			[7:0] in_data244;
reg			[7:0] in_data245;
reg			[7:0] in_data246;
reg			[7:0] in_data247;
reg			[7:0] in_data248;
reg			[7:0] in_data249;
reg			[7:0] in_data250;
reg			[7:0] in_data251;
reg			[7:0] in_data252;
reg			[7:0] in_data253;
reg			[7:0] in_data254;
reg			[7:0] in_data255;






/*
 * Store input into memory
 */
reg			[8:0] input_index;
reg				  in_valid_flag; //so that calculation of bubble sort can start right after in_valid is low
reg				  bubble_start_flag; //indicates the start of bubble sort (combinational)
always @(posedge clk) begin
	if (!rst_n) begin
		input_index <= 'd0;
		in_valid_flag <= 1'b0;
		bubble_start_flag <= 1'b0;
		in_data0 <= 'd0;
		in_data1 <= 'd0;
		in_data2 <= 'd0;
		in_data3 <= 'd0;
		in_data4 <= 'd0;
		in_data5 <= 'd0;
		in_data6 <= 'd0;
		in_data7 <= 'd0;
		in_data8 <= 'd0;
		in_data9 <= 'd0;
		in_data10 <= 'd0;
		in_data11 <= 'd0;
		in_data12 <= 'd0;
		in_data13 <= 'd0;
		in_data14 <= 'd0;
		in_data15 <= 'd0;
		in_data16 <= 'd0;
		in_data17 <= 'd0;
		in_data18 <= 'd0;
		in_data19 <= 'd0;
		in_data20 <= 'd0;
		in_data21 <= 'd0;
		in_data22 <= 'd0;
		in_data23 <= 'd0;
		in_data24 <= 'd0;
		in_data25 <= 'd0;
		in_data26 <= 'd0;
		in_data27 <= 'd0;
		in_data28 <= 'd0;
		in_data29 <= 'd0;
		in_data30 <= 'd0;
		in_data31 <= 'd0;
		in_data32 <= 'd0;
		in_data33 <= 'd0;
		in_data34 <= 'd0;
		in_data35 <= 'd0;
		in_data36 <= 'd0;
		in_data37 <= 'd0;
		in_data38 <= 'd0;
		in_data39 <= 'd0;
		in_data40 <= 'd0;
		in_data41 <= 'd0;
		in_data42 <= 'd0;
		in_data43 <= 'd0;
		in_data44 <= 'd0;
		in_data45 <= 'd0;
		in_data46 <= 'd0;
		in_data47 <= 'd0;
		in_data48 <= 'd0;
		in_data49 <= 'd0;
		in_data50 <= 'd0;
		in_data51 <= 'd0;
		in_data52 <= 'd0;
		in_data53 <= 'd0;
		in_data54 <= 'd0;
		in_data55 <= 'd0;
		in_data56 <= 'd0;
		in_data57 <= 'd0;
		in_data58 <= 'd0;
		in_data59 <= 'd0;
		in_data60 <= 'd0;
		in_data61 <= 'd0;
		in_data62 <= 'd0;
		in_data63 <= 'd0;
		in_data64 <= 'd0;
		in_data65 <= 'd0;
		in_data66 <= 'd0;
		in_data67 <= 'd0;
		in_data68 <= 'd0;
		in_data69 <= 'd0;
		in_data70 <= 'd0;
		in_data71 <= 'd0;
		in_data72 <= 'd0;
		in_data73 <= 'd0;
		in_data74 <= 'd0;
		in_data75 <= 'd0;
		in_data76 <= 'd0;
		in_data77 <= 'd0;
		in_data78 <= 'd0;
		in_data79 <= 'd0;
		in_data80 <= 'd0;
		in_data81 <= 'd0;
		in_data82 <= 'd0;
		in_data83 <= 'd0;
		in_data84 <= 'd0;
		in_data85 <= 'd0;
		in_data86 <= 'd0;
		in_data87 <= 'd0;
		in_data88 <= 'd0;
		in_data89 <= 'd0;
		in_data90 <= 'd0;
		in_data91 <= 'd0;
		in_data92 <= 'd0;
		in_data93 <= 'd0;
		in_data94 <= 'd0;
		in_data95 <= 'd0;
		in_data96 <= 'd0;
		in_data97 <= 'd0;
		in_data98 <= 'd0;
		in_data99 <= 'd0;
		in_data100 <= 'd0;
		in_data101 <= 'd0;
		in_data102 <= 'd0;
		in_data103 <= 'd0;
		in_data104 <= 'd0;
		in_data105 <= 'd0;
		in_data106 <= 'd0;
		in_data107 <= 'd0;
		in_data108 <= 'd0;
		in_data109 <= 'd0;
		in_data110 <= 'd0;
		in_data111 <= 'd0;
		in_data112 <= 'd0;
		in_data113 <= 'd0;
		in_data114 <= 'd0;
		in_data115 <= 'd0;
		in_data116 <= 'd0;
		in_data117 <= 'd0;
		in_data118 <= 'd0;
		in_data119 <= 'd0;
		in_data120 <= 'd0;
		in_data121 <= 'd0;
		in_data122 <= 'd0;
		in_data123 <= 'd0;
		in_data124 <= 'd0;
		in_data125 <= 'd0;
		in_data126 <= 'd0;
		in_data127 <= 'd0;
		in_data128 <= 'd0;
		in_data129 <= 'd0;
		in_data130 <= 'd0;
		in_data131 <= 'd0;
		in_data132 <= 'd0;
		in_data133 <= 'd0;
		in_data134 <= 'd0;
		in_data135 <= 'd0;
		in_data136 <= 'd0;
		in_data137 <= 'd0;
		in_data138 <= 'd0;
		in_data139 <= 'd0;
		in_data140 <= 'd0;
		in_data141 <= 'd0;
		in_data142 <= 'd0;
		in_data143 <= 'd0;
		in_data144 <= 'd0;
		in_data145 <= 'd0;
		in_data146 <= 'd0;
		in_data147 <= 'd0;
		in_data148 <= 'd0;
		in_data149 <= 'd0;
		in_data150 <= 'd0;
		in_data151 <= 'd0;
		in_data152 <= 'd0;
		in_data153 <= 'd0;
		in_data154 <= 'd0;
		in_data155 <= 'd0;
		in_data156 <= 'd0;
		in_data157 <= 'd0;
		in_data158 <= 'd0;
		in_data159 <= 'd0;
		in_data160 <= 'd0;
		in_data161 <= 'd0;
		in_data162 <= 'd0;
		in_data163 <= 'd0;
		in_data164 <= 'd0;
		in_data165 <= 'd0;
		in_data166 <= 'd0;
		in_data167 <= 'd0;
		in_data168 <= 'd0;
		in_data169 <= 'd0;
		in_data170 <= 'd0;
		in_data171 <= 'd0;
		in_data172 <= 'd0;
		in_data173 <= 'd0;
		in_data174 <= 'd0;
		in_data175 <= 'd0;
		in_data176 <= 'd0;
		in_data177 <= 'd0;
		in_data178 <= 'd0;
		in_data179 <= 'd0;
		in_data180 <= 'd0;
		in_data181 <= 'd0;
		in_data182 <= 'd0;
		in_data183 <= 'd0;
		in_data184 <= 'd0;
		in_data185 <= 'd0;
		in_data186 <= 'd0;
		in_data187 <= 'd0;
		in_data188 <= 'd0;
		in_data189 <= 'd0;
		in_data190 <= 'd0;
		in_data191 <= 'd0;
		in_data192 <= 'd0;
		in_data193 <= 'd0;
		in_data194 <= 'd0;
		in_data195 <= 'd0;
		in_data196 <= 'd0;
		in_data197 <= 'd0;
		in_data198 <= 'd0;
		in_data199 <= 'd0;
		in_data200 <= 'd0;
		in_data201 <= 'd0;
		in_data202 <= 'd0;
		in_data203 <= 'd0;
		in_data204 <= 'd0;
		in_data205 <= 'd0;
		in_data206 <= 'd0;
		in_data207 <= 'd0;
		in_data208 <= 'd0;
		in_data209 <= 'd0;
		in_data210 <= 'd0;
		in_data211 <= 'd0;
		in_data212 <= 'd0;
		in_data213 <= 'd0;
		in_data214 <= 'd0;
		in_data215 <= 'd0;
		in_data216 <= 'd0;
		in_data217 <= 'd0;
		in_data218 <= 'd0;
		in_data219 <= 'd0;
		in_data220 <= 'd0;
		in_data221 <= 'd0;
		in_data222 <= 'd0;
		in_data223 <= 'd0;
		in_data224 <= 'd0;
		in_data225 <= 'd0;
		in_data226 <= 'd0;
		in_data227 <= 'd0;
		in_data228 <= 'd0;
		in_data229 <= 'd0;
		in_data230 <= 'd0;
		in_data231 <= 'd0;
		in_data232 <= 'd0;
		in_data233 <= 'd0;
		in_data234 <= 'd0;
		in_data235 <= 'd0;
		in_data236 <= 'd0;
		in_data237 <= 'd0;
		in_data238 <= 'd0;
		in_data239 <= 'd0;
		in_data240 <= 'd0;
		in_data241 <= 'd0;
		in_data242 <= 'd0;
		in_data243 <= 'd0;
		in_data244 <= 'd0;
		in_data245 <= 'd0;
		in_data246 <= 'd0;
		in_data247 <= 'd0;
		in_data248 <= 'd0;
		in_data249 <= 'd0;
		in_data250 <= 'd0;
		in_data251 <= 'd0;
		in_data252 <= 'd0;
		in_data253 <= 'd0;
		in_data254 <= 'd0;
		in_data255 <= 'd0;
	end
	else begin
		if(in_valid) begin
			in_valid_flag <= 1'b1;
			input_index <= input_index + 1'b1;

			case(input_index)
				'd0: in_data0 <= in_data;
				'd1: in_data1 <= in_data;
				'd2: in_data2 <= in_data;
				'd3: in_data3 <= in_data;
				'd4: in_data4 <= in_data;
				'd5: in_data5 <= in_data;
				'd6: in_data6 <= in_data;
				'd7: in_data7 <= in_data;
				'd8: in_data8 <= in_data;
				'd9: in_data9 <= in_data;
				'd10: in_data10 <= in_data;
				'd11: in_data11 <= in_data;
				'd12: in_data12 <= in_data;
				'd13: in_data13 <= in_data;
				'd14: in_data14 <= in_data;
				'd15: in_data15 <= in_data;
				'd16: in_data16 <= in_data;
				'd17: in_data17 <= in_data;
				'd18: in_data18 <= in_data;
				'd19: in_data19 <= in_data;
				'd20: in_data20 <= in_data;
				'd21: in_data21 <= in_data;
				'd22: in_data22 <= in_data;
				'd23: in_data23 <= in_data;
				'd24: in_data24 <= in_data;
				'd25: in_data25 <= in_data;
				'd26: in_data26 <= in_data;
				'd27: in_data27 <= in_data;
				'd28: in_data28 <= in_data;
				'd29: in_data29 <= in_data;
				'd30: in_data30 <= in_data;
				'd31: in_data31 <= in_data;
				'd32: in_data32 <= in_data;
				'd33: in_data33 <= in_data;
				'd34: in_data34 <= in_data;
				'd35: in_data35 <= in_data;
				'd36: in_data36 <= in_data;
				'd37: in_data37 <= in_data;
				'd38: in_data38 <= in_data;
				'd39: in_data39 <= in_data;
				'd40: in_data40 <= in_data;
				'd41: in_data41 <= in_data;
				'd42: in_data42 <= in_data;
				'd43: in_data43 <= in_data;
				'd44: in_data44 <= in_data;
				'd45: in_data45 <= in_data;
				'd46: in_data46 <= in_data;
				'd47: in_data47 <= in_data;
				'd48: in_data48 <= in_data;
				'd49: in_data49 <= in_data;
				'd50: in_data50 <= in_data;
				'd51: in_data51 <= in_data;
				'd52: in_data52 <= in_data;
				'd53: in_data53 <= in_data;
				'd54: in_data54 <= in_data;
				'd55: in_data55 <= in_data;
				'd56: in_data56 <= in_data;
				'd57: in_data57 <= in_data;
				'd58: in_data58 <= in_data;
				'd59: in_data59 <= in_data;
				'd60: in_data60 <= in_data;
				'd61: in_data61 <= in_data;
				'd62: in_data62 <= in_data;
				'd63: in_data63 <= in_data;
				'd64: in_data64 <= in_data;
				'd65: in_data65 <= in_data;
				'd66: in_data66 <= in_data;
				'd67: in_data67 <= in_data;
				'd68: in_data68 <= in_data;
				'd69: in_data69 <= in_data;
				'd70: in_data70 <= in_data;
				'd71: in_data71 <= in_data;
				'd72: in_data72 <= in_data;
				'd73: in_data73 <= in_data;
				'd74: in_data74 <= in_data;
				'd75: in_data75 <= in_data;
				'd76: in_data76 <= in_data;
				'd77: in_data77 <= in_data;
				'd78: in_data78 <= in_data;
				'd79: in_data79 <= in_data;
				'd80: in_data80 <= in_data;
				'd81: in_data81 <= in_data;
				'd82: in_data82 <= in_data;
				'd83: in_data83 <= in_data;
				'd84: in_data84 <= in_data;
				'd85: in_data85 <= in_data;
				'd86: in_data86 <= in_data;
				'd87: in_data87 <= in_data;
				'd88: in_data88 <= in_data;
				'd89: in_data89 <= in_data;
				'd90: in_data90 <= in_data;
				'd91: in_data91 <= in_data;
				'd92: in_data92 <= in_data;
				'd93: in_data93 <= in_data;
				'd94: in_data94 <= in_data;
				'd95: in_data95 <= in_data;
				'd96: in_data96 <= in_data;
				'd97: in_data97 <= in_data;
				'd98: in_data98 <= in_data;
				'd99: in_data99 <= in_data;
				'd100: in_data100 <= in_data;
				'd101: in_data101 <= in_data;
				'd102: in_data102 <= in_data;
				'd103: in_data103 <= in_data;
				'd104: in_data104 <= in_data;
				'd105: in_data105 <= in_data;
				'd106: in_data106 <= in_data;
				'd107: in_data107 <= in_data;
				'd108: in_data108 <= in_data;
				'd109: in_data109 <= in_data;
				'd110: in_data110 <= in_data;
				'd111: in_data111 <= in_data;
				'd112: in_data112 <= in_data;
				'd113: in_data113 <= in_data;
				'd114: in_data114 <= in_data;
				'd115: in_data115 <= in_data;
				'd116: in_data116 <= in_data;
				'd117: in_data117 <= in_data;
				'd118: in_data118 <= in_data;
				'd119: in_data119 <= in_data;
				'd120: in_data120 <= in_data;
				'd121: in_data121 <= in_data;
				'd122: in_data122 <= in_data;
				'd123: in_data123 <= in_data;
				'd124: in_data124 <= in_data;
				'd125: in_data125 <= in_data;
				'd126: in_data126 <= in_data;
				'd127: in_data127 <= in_data;
				'd128: in_data128 <= in_data;
				'd129: in_data129 <= in_data;
				'd130: in_data130 <= in_data;
				'd131: in_data131 <= in_data;
				'd132: in_data132 <= in_data;
				'd133: in_data133 <= in_data;
				'd134: in_data134 <= in_data;
				'd135: in_data135 <= in_data;
				'd136: in_data136 <= in_data;
				'd137: in_data137 <= in_data;
				'd138: in_data138 <= in_data;
				'd139: in_data139 <= in_data;
				'd140: in_data140 <= in_data;
				'd141: in_data141 <= in_data;
				'd142: in_data142 <= in_data;
				'd143: in_data143 <= in_data;
				'd144: in_data144 <= in_data;
				'd145: in_data145 <= in_data;
				'd146: in_data146 <= in_data;
				'd147: in_data147 <= in_data;
				'd148: in_data148 <= in_data;
				'd149: in_data149 <= in_data;
				'd150: in_data150 <= in_data;
				'd151: in_data151 <= in_data;
				'd152: in_data152 <= in_data;
				'd153: in_data153 <= in_data;
				'd154: in_data154 <= in_data;
				'd155: in_data155 <= in_data;
				'd156: in_data156 <= in_data;
				'd157: in_data157 <= in_data;
				'd158: in_data158 <= in_data;
				'd159: in_data159 <= in_data;
				'd160: in_data160 <= in_data;
				'd161: in_data161 <= in_data;
				'd162: in_data162 <= in_data;
				'd163: in_data163 <= in_data;
				'd164: in_data164 <= in_data;
				'd165: in_data165 <= in_data;
				'd166: in_data166 <= in_data;
				'd167: in_data167 <= in_data;
				'd168: in_data168 <= in_data;
				'd169: in_data169 <= in_data;
				'd170: in_data170 <= in_data;
				'd171: in_data171 <= in_data;
				'd172: in_data172 <= in_data;
				'd173: in_data173 <= in_data;
				'd174: in_data174 <= in_data;
				'd175: in_data175 <= in_data;
				'd176: in_data176 <= in_data;
				'd177: in_data177 <= in_data;
				'd178: in_data178 <= in_data;
				'd179: in_data179 <= in_data;
				'd180: in_data180 <= in_data;
				'd181: in_data181 <= in_data;
				'd182: in_data182 <= in_data;
				'd183: in_data183 <= in_data;
				'd184: in_data184 <= in_data;
				'd185: in_data185 <= in_data;
				'd186: in_data186 <= in_data;
				'd187: in_data187 <= in_data;
				'd188: in_data188 <= in_data;
				'd189: in_data189 <= in_data;
				'd190: in_data190 <= in_data;
				'd191: in_data191 <= in_data;
				'd192: in_data192 <= in_data;
				'd193: in_data193 <= in_data;
				'd194: in_data194 <= in_data;
				'd195: in_data195 <= in_data;
				'd196: in_data196 <= in_data;
				'd197: in_data197 <= in_data;
				'd198: in_data198 <= in_data;
				'd199: in_data199 <= in_data;
				'd200: in_data200 <= in_data;
				'd201: in_data201 <= in_data;
				'd202: in_data202 <= in_data;
				'd203: in_data203 <= in_data;
				'd204: in_data204 <= in_data;
				'd205: in_data205 <= in_data;
				'd206: in_data206 <= in_data;
				'd207: in_data207 <= in_data;
				'd208: in_data208 <= in_data;
				'd209: in_data209 <= in_data;
				'd210: in_data210 <= in_data;
				'd211: in_data211 <= in_data;
				'd212: in_data212 <= in_data;
				'd213: in_data213 <= in_data;
				'd214: in_data214 <= in_data;
				'd215: in_data215 <= in_data;
				'd216: in_data216 <= in_data;
				'd217: in_data217 <= in_data;
				'd218: in_data218 <= in_data;
				'd219: in_data219 <= in_data;
				'd220: in_data220 <= in_data;
				'd221: in_data221 <= in_data;
				'd222: in_data222 <= in_data;
				'd223: in_data223 <= in_data;
				'd224: in_data224 <= in_data;
				'd225: in_data225 <= in_data;
				'd226: in_data226 <= in_data;
				'd227: in_data227 <= in_data;
				'd228: in_data228 <= in_data;
				'd229: in_data229 <= in_data;
				'd230: in_data230 <= in_data;
				'd231: in_data231 <= in_data;
				'd232: in_data232 <= in_data;
				'd233: in_data233 <= in_data;
				'd234: in_data234 <= in_data;
				'd235: in_data235 <= in_data;
				'd236: in_data236 <= in_data;
				'd237: in_data237 <= in_data;
				'd238: in_data238 <= in_data;
				'd239: in_data239 <= in_data;
				'd240: in_data240 <= in_data;
				'd241: in_data241 <= in_data;
				'd242: in_data242 <= in_data;
				'd243: in_data243 <= in_data;
				'd244: in_data244 <= in_data;
				'd245: in_data245 <= in_data;
				'd246: in_data246 <= in_data;
				'd247: in_data247 <= in_data;
				'd248: in_data248 <= in_data;
				'd249: in_data249 <= in_data;
				'd250: in_data250 <= in_data;
				'd251: in_data251 <= in_data;
				'd252: in_data252 <= in_data;
				'd253: in_data253 <= in_data;
				'd254: in_data254 <= in_data;
				'd255: in_data255 <= in_data;
			endcase
		end
		else begin//!in_valid
			if(dump_out_flag) begin
				input_index <= 'd0;
				bubble_start_flag <= 1'b0;
				in_valid_flag <= 1'b0;

				//Clear Input Datas
				in_data0 <= 'd0;
				in_data1 <= 'd0;
				in_data2 <= 'd0;
				in_data3 <= 'd0;
				in_data4 <= 'd0;
				in_data5 <= 'd0;
				in_data6 <= 'd0;
				in_data7 <= 'd0;
				in_data8 <= 'd0;
				in_data9 <= 'd0;
				in_data10 <= 'd0;
				in_data11 <= 'd0;
				in_data12 <= 'd0;
				in_data13 <= 'd0;
				in_data14 <= 'd0;
				in_data15 <= 'd0;
				in_data16 <= 'd0;
				in_data17 <= 'd0;
				in_data18 <= 'd0;
				in_data19 <= 'd0;
				in_data20 <= 'd0;
				in_data21 <= 'd0;
				in_data22 <= 'd0;
				in_data23 <= 'd0;
				in_data24 <= 'd0;
				in_data25 <= 'd0;
				in_data26 <= 'd0;
				in_data27 <= 'd0;
				in_data28 <= 'd0;
				in_data29 <= 'd0;
				in_data30 <= 'd0;
				in_data31 <= 'd0;
				in_data32 <= 'd0;
				in_data33 <= 'd0;
				in_data34 <= 'd0;
				in_data35 <= 'd0;
				in_data36 <= 'd0;
				in_data37 <= 'd0;
				in_data38 <= 'd0;
				in_data39 <= 'd0;
				in_data40 <= 'd0;
				in_data41 <= 'd0;
				in_data42 <= 'd0;
				in_data43 <= 'd0;
				in_data44 <= 'd0;
				in_data45 <= 'd0;
				in_data46 <= 'd0;
				in_data47 <= 'd0;
				in_data48 <= 'd0;
				in_data49 <= 'd0;
				in_data50 <= 'd0;
				in_data51 <= 'd0;
				in_data52 <= 'd0;
				in_data53 <= 'd0;
				in_data54 <= 'd0;
				in_data55 <= 'd0;
				in_data56 <= 'd0;
				in_data57 <= 'd0;
				in_data58 <= 'd0;
				in_data59 <= 'd0;
				in_data60 <= 'd0;
				in_data61 <= 'd0;
				in_data62 <= 'd0;
				in_data63 <= 'd0;
				in_data64 <= 'd0;
				in_data65 <= 'd0;
				in_data66 <= 'd0;
				in_data67 <= 'd0;
				in_data68 <= 'd0;
				in_data69 <= 'd0;
				in_data70 <= 'd0;
				in_data71 <= 'd0;
				in_data72 <= 'd0;
				in_data73 <= 'd0;
				in_data74 <= 'd0;
				in_data75 <= 'd0;
				in_data76 <= 'd0;
				in_data77 <= 'd0;
				in_data78 <= 'd0;
				in_data79 <= 'd0;
				in_data80 <= 'd0;
				in_data81 <= 'd0;
				in_data82 <= 'd0;
				in_data83 <= 'd0;
				in_data84 <= 'd0;
				in_data85 <= 'd0;
				in_data86 <= 'd0;
				in_data87 <= 'd0;
				in_data88 <= 'd0;
				in_data89 <= 'd0;
				in_data90 <= 'd0;
				in_data91 <= 'd0;
				in_data92 <= 'd0;
				in_data93 <= 'd0;
				in_data94 <= 'd0;
				in_data95 <= 'd0;
				in_data96 <= 'd0;
				in_data97 <= 'd0;
				in_data98 <= 'd0;
				in_data99 <= 'd0;
				in_data100 <= 'd0;
				in_data101 <= 'd0;
				in_data102 <= 'd0;
				in_data103 <= 'd0;
				in_data104 <= 'd0;
				in_data105 <= 'd0;
				in_data106 <= 'd0;
				in_data107 <= 'd0;
				in_data108 <= 'd0;
				in_data109 <= 'd0;
				in_data110 <= 'd0;
				in_data111 <= 'd0;
				in_data112 <= 'd0;
				in_data113 <= 'd0;
				in_data114 <= 'd0;
				in_data115 <= 'd0;
				in_data116 <= 'd0;
				in_data117 <= 'd0;
				in_data118 <= 'd0;
				in_data119 <= 'd0;
				in_data120 <= 'd0;
				in_data121 <= 'd0;
				in_data122 <= 'd0;
				in_data123 <= 'd0;
				in_data124 <= 'd0;
				in_data125 <= 'd0;
				in_data126 <= 'd0;
				in_data127 <= 'd0;
				in_data128 <= 'd0;
				in_data129 <= 'd0;
				in_data130 <= 'd0;
				in_data131 <= 'd0;
				in_data132 <= 'd0;
				in_data133 <= 'd0;
				in_data134 <= 'd0;
				in_data135 <= 'd0;
				in_data136 <= 'd0;
				in_data137 <= 'd0;
				in_data138 <= 'd0;
				in_data139 <= 'd0;
				in_data140 <= 'd0;
				in_data141 <= 'd0;
				in_data142 <= 'd0;
				in_data143 <= 'd0;
				in_data144 <= 'd0;
				in_data145 <= 'd0;
				in_data146 <= 'd0;
				in_data147 <= 'd0;
				in_data148 <= 'd0;
				in_data149 <= 'd0;
				in_data150 <= 'd0;
				in_data151 <= 'd0;
				in_data152 <= 'd0;
				in_data153 <= 'd0;
				in_data154 <= 'd0;
				in_data155 <= 'd0;
				in_data156 <= 'd0;
				in_data157 <= 'd0;
				in_data158 <= 'd0;
				in_data159 <= 'd0;
				in_data160 <= 'd0;
				in_data161 <= 'd0;
				in_data162 <= 'd0;
				in_data163 <= 'd0;
				in_data164 <= 'd0;
				in_data165 <= 'd0;
				in_data166 <= 'd0;
				in_data167 <= 'd0;
				in_data168 <= 'd0;
				in_data169 <= 'd0;
				in_data170 <= 'd0;
				in_data171 <= 'd0;
				in_data172 <= 'd0;
				in_data173 <= 'd0;
				in_data174 <= 'd0;
				in_data175 <= 'd0;
				in_data176 <= 'd0;
				in_data177 <= 'd0;
				in_data178 <= 'd0;
				in_data179 <= 'd0;
				in_data180 <= 'd0;
				in_data181 <= 'd0;
				in_data182 <= 'd0;
				in_data183 <= 'd0;
				in_data184 <= 'd0;
				in_data185 <= 'd0;
				in_data186 <= 'd0;
				in_data187 <= 'd0;
				in_data188 <= 'd0;
				in_data189 <= 'd0;
				in_data190 <= 'd0;
				in_data191 <= 'd0;
				in_data192 <= 'd0;
				in_data193 <= 'd0;
				in_data194 <= 'd0;
				in_data195 <= 'd0;
				in_data196 <= 'd0;
				in_data197 <= 'd0;
				in_data198 <= 'd0;
				in_data199 <= 'd0;
				in_data200 <= 'd0;
				in_data201 <= 'd0;
				in_data202 <= 'd0;
				in_data203 <= 'd0;
				in_data204 <= 'd0;
				in_data205 <= 'd0;
				in_data206 <= 'd0;
				in_data207 <= 'd0;
				in_data208 <= 'd0;
				in_data209 <= 'd0;
				in_data210 <= 'd0;
				in_data211 <= 'd0;
				in_data212 <= 'd0;
				in_data213 <= 'd0;
				in_data214 <= 'd0;
				in_data215 <= 'd0;
				in_data216 <= 'd0;
				in_data217 <= 'd0;
				in_data218 <= 'd0;
				in_data219 <= 'd0;
				in_data220 <= 'd0;
				in_data221 <= 'd0;
				in_data222 <= 'd0;
				in_data223 <= 'd0;
				in_data224 <= 'd0;
				in_data225 <= 'd0;
				in_data226 <= 'd0;
				in_data227 <= 'd0;
				in_data228 <= 'd0;
				in_data229 <= 'd0;
				in_data230 <= 'd0;
				in_data231 <= 'd0;
				in_data232 <= 'd0;
				in_data233 <= 'd0;
				in_data234 <= 'd0;
				in_data235 <= 'd0;
				in_data236 <= 'd0;
				in_data237 <= 'd0;
				in_data238 <= 'd0;
				in_data239 <= 'd0;
				in_data240 <= 'd0;
				in_data241 <= 'd0;
				in_data242 <= 'd0;
				in_data243 <= 'd0;
				in_data244 <= 'd0;
				in_data245 <= 'd0;
				in_data246 <= 'd0;
				in_data247 <= 'd0;
				in_data248 <= 'd0;
				in_data249 <= 'd0;
				in_data250 <= 'd0;
				in_data251 <= 'd0;
				in_data252 <= 'd0;
				in_data253 <= 'd0;
				in_data254 <= 'd0;
				in_data255 <= 'd0;
			end
			else if(in_valid_flag) begin
				bubble_start_flag <= 1'b1;
			end
			else begin
				bubble_start_flag <= 1'b0;
			end
		end
	end
end



/*
 * Bubble Sort
 * -------------
 * - Break into ODD and EVEN parts
 * - INDEX of OUTER LOOP set to # of INPUTS (for now)
 */

reg				[8:0] outer_loop;
always @(posedge clk) begin
	if (!rst_n) begin
		outer_loop <= 'd0;	
	end
	else if (bubble_start_flag) begin
		if(outer_loop < input_index) begin
			outer_loop <= outer_loop + 1'b1;
		end
		else if(dump_out_flag) begin//finish dumping outputs
			outer_loop <= 'd0;
		end
		else begin
			outer_loop <= outer_loop;
		end
	end
end





/*
 * Dump Output
 */
 reg			[8:0] output_index;
always @(posedge clk) begin
	if (!rst_n) begin
		output_index <= 'd0;		
	end
	else if (dump_out_flag) begin
		dump_out_flag <= 1'b0;
		output_index <= 'd0;
	end
	else if (outer_loop == input_index) begin//sorted for outer_loop # of times
		if (output_index < input_index) begin
			output_index <= output_index + 1'b1;
			out_valid <= 1'b1;
			case(output_index)
				'd0: out_data <= in_data0;
				'd1: out_data <= in_data1;
				'd2: out_data <= in_data2;
				'd3: out_data <= in_data3;
				'd4: out_data <= in_data4;
				'd5: out_data <= in_data5;
				'd6: out_data <= in_data6;
				'd7: out_data <= in_data7;
				'd8: out_data <= in_data8;
				'd9: out_data <= in_data9;
				'd10: out_data <= in_data10;
				'd11: out_data <= in_data11;
				'd12: out_data <= in_data12;
				'd13: out_data <= in_data13;
				'd14: out_data <= in_data14;
				'd15: out_data <= in_data15;
				'd16: out_data <= in_data16;
				'd17: out_data <= in_data17;
				'd18: out_data <= in_data18;
				'd19: out_data <= in_data19;
				'd20: out_data <= in_data20;
				'd21: out_data <= in_data21;
				'd22: out_data <= in_data22;
				'd23: out_data <= in_data23;
				'd24: out_data <= in_data24;
				'd25: out_data <= in_data25;
				'd26: out_data <= in_data26;
				'd27: out_data <= in_data27;
				'd28: out_data <= in_data28;
				'd29: out_data <= in_data29;
				'd30: out_data <= in_data30;
				'd31: out_data <= in_data31;
				'd32: out_data <= in_data32;
				'd33: out_data <= in_data33;
				'd34: out_data <= in_data34;
				'd35: out_data <= in_data35;
				'd36: out_data <= in_data36;
				'd37: out_data <= in_data37;
				'd38: out_data <= in_data38;
				'd39: out_data <= in_data39;
				'd40: out_data <= in_data40;
				'd41: out_data <= in_data41;
				'd42: out_data <= in_data42;
				'd43: out_data <= in_data43;
				'd44: out_data <= in_data44;
				'd45: out_data <= in_data45;
				'd46: out_data <= in_data46;
				'd47: out_data <= in_data47;
				'd48: out_data <= in_data48;
				'd49: out_data <= in_data49;
				'd50: out_data <= in_data50;
				'd51: out_data <= in_data51;
				'd52: out_data <= in_data52;
				'd53: out_data <= in_data53;
				'd54: out_data <= in_data54;
				'd55: out_data <= in_data55;
				'd56: out_data <= in_data56;
				'd57: out_data <= in_data57;
				'd58: out_data <= in_data58;
				'd59: out_data <= in_data59;
				'd60: out_data <= in_data60;
				'd61: out_data <= in_data61;
				'd62: out_data <= in_data62;
				'd63: out_data <= in_data63;
				'd64: out_data <= in_data64;
				'd65: out_data <= in_data65;
				'd66: out_data <= in_data66;
				'd67: out_data <= in_data67;
				'd68: out_data <= in_data68;
				'd69: out_data <= in_data69;
				'd70: out_data <= in_data70;
				'd71: out_data <= in_data71;
				'd72: out_data <= in_data72;
				'd73: out_data <= in_data73;
				'd74: out_data <= in_data74;
				'd75: out_data <= in_data75;
				'd76: out_data <= in_data76;
				'd77: out_data <= in_data77;
				'd78: out_data <= in_data78;
				'd79: out_data <= in_data79;
				'd80: out_data <= in_data80;
				'd81: out_data <= in_data81;
				'd82: out_data <= in_data82;
				'd83: out_data <= in_data83;
				'd84: out_data <= in_data84;
				'd85: out_data <= in_data85;
				'd86: out_data <= in_data86;
				'd87: out_data <= in_data87;
				'd88: out_data <= in_data88;
				'd89: out_data <= in_data89;
				'd90: out_data <= in_data90;
				'd91: out_data <= in_data91;
				'd92: out_data <= in_data92;
				'd93: out_data <= in_data93;
				'd94: out_data <= in_data94;
				'd95: out_data <= in_data95;
				'd96: out_data <= in_data96;
				'd97: out_data <= in_data97;
				'd98: out_data <= in_data98;
				'd99: out_data <= in_data99;
				'd100: out_data <= in_data100;
				'd101: out_data <= in_data101;
				'd102: out_data <= in_data102;
				'd103: out_data <= in_data103;
				'd104: out_data <= in_data104;
				'd105: out_data <= in_data105;
				'd106: out_data <= in_data106;
				'd107: out_data <= in_data107;
				'd108: out_data <= in_data108;
				'd109: out_data <= in_data109;
				'd110: out_data <= in_data110;
				'd111: out_data <= in_data111;
				'd112: out_data <= in_data112;
				'd113: out_data <= in_data113;
				'd114: out_data <= in_data114;
				'd115: out_data <= in_data115;
				'd116: out_data <= in_data116;
				'd117: out_data <= in_data117;
				'd118: out_data <= in_data118;
				'd119: out_data <= in_data119;
				'd120: out_data <= in_data120;
				'd121: out_data <= in_data121;
				'd122: out_data <= in_data122;
				'd123: out_data <= in_data123;
				'd124: out_data <= in_data124;
				'd125: out_data <= in_data125;
				'd126: out_data <= in_data126;
				'd127: out_data <= in_data127;
				'd128: out_data <= in_data128;
				'd129: out_data <= in_data129;
				'd130: out_data <= in_data130;
				'd131: out_data <= in_data131;
				'd132: out_data <= in_data132;
				'd133: out_data <= in_data133;
				'd134: out_data <= in_data134;
				'd135: out_data <= in_data135;
				'd136: out_data <= in_data136;
				'd137: out_data <= in_data137;
				'd138: out_data <= in_data138;
				'd139: out_data <= in_data139;
				'd140: out_data <= in_data140;
				'd141: out_data <= in_data141;
				'd142: out_data <= in_data142;
				'd143: out_data <= in_data143;
				'd144: out_data <= in_data144;
				'd145: out_data <= in_data145;
				'd146: out_data <= in_data146;
				'd147: out_data <= in_data147;
				'd148: out_data <= in_data148;
				'd149: out_data <= in_data149;
				'd150: out_data <= in_data150;
				'd151: out_data <= in_data151;
				'd152: out_data <= in_data152;
				'd153: out_data <= in_data153;
				'd154: out_data <= in_data154;
				'd155: out_data <= in_data155;
				'd156: out_data <= in_data156;
				'd157: out_data <= in_data157;
				'd158: out_data <= in_data158;
				'd159: out_data <= in_data159;
				'd160: out_data <= in_data160;
				'd161: out_data <= in_data161;
				'd162: out_data <= in_data162;
				'd163: out_data <= in_data163;
				'd164: out_data <= in_data164;
				'd165: out_data <= in_data165;
				'd166: out_data <= in_data166;
				'd167: out_data <= in_data167;
				'd168: out_data <= in_data168;
				'd169: out_data <= in_data169;
				'd170: out_data <= in_data170;
				'd171: out_data <= in_data171;
				'd172: out_data <= in_data172;
				'd173: out_data <= in_data173;
				'd174: out_data <= in_data174;
				'd175: out_data <= in_data175;
				'd176: out_data <= in_data176;
				'd177: out_data <= in_data177;
				'd178: out_data <= in_data178;
				'd179: out_data <= in_data179;
				'd180: out_data <= in_data180;
				'd181: out_data <= in_data181;
				'd182: out_data <= in_data182;
				'd183: out_data <= in_data183;
				'd184: out_data <= in_data184;
				'd185: out_data <= in_data185;
				'd186: out_data <= in_data186;
				'd187: out_data <= in_data187;
				'd188: out_data <= in_data188;
				'd189: out_data <= in_data189;
				'd190: out_data <= in_data190;
				'd191: out_data <= in_data191;
				'd192: out_data <= in_data192;
				'd193: out_data <= in_data193;
				'd194: out_data <= in_data194;
				'd195: out_data <= in_data195;
				'd196: out_data <= in_data196;
				'd197: out_data <= in_data197;
				'd198: out_data <= in_data198;
				'd199: out_data <= in_data199;
				'd200: out_data <= in_data200;
				'd201: out_data <= in_data201;
				'd202: out_data <= in_data202;
				'd203: out_data <= in_data203;
				'd204: out_data <= in_data204;
				'd205: out_data <= in_data205;
				'd206: out_data <= in_data206;
				'd207: out_data <= in_data207;
				'd208: out_data <= in_data208;
				'd209: out_data <= in_data209;
				'd210: out_data <= in_data210;
				'd211: out_data <= in_data211;
				'd212: out_data <= in_data212;
				'd213: out_data <= in_data213;
				'd214: out_data <= in_data214;
				'd215: out_data <= in_data215;
				'd216: out_data <= in_data216;
				'd217: out_data <= in_data217;
				'd218: out_data <= in_data218;
				'd219: out_data <= in_data219;
				'd220: out_data <= in_data220;
				'd221: out_data <= in_data221;
				'd222: out_data <= in_data222;
				'd223: out_data <= in_data223;
				'd224: out_data <= in_data224;
				'd225: out_data <= in_data225;
				'd226: out_data <= in_data226;
				'd227: out_data <= in_data227;
				'd228: out_data <= in_data228;
				'd229: out_data <= in_data229;
				'd230: out_data <= in_data230;
				'd231: out_data <= in_data231;
				'd232: out_data <= in_data232;
				'd233: out_data <= in_data233;
				'd234: out_data <= in_data234;
				'd235: out_data <= in_data235;
				'd236: out_data <= in_data236;
				'd237: out_data <= in_data237;
				'd238: out_data <= in_data238;
				'd239: out_data <= in_data239;
				'd240: out_data <= in_data240;
				'd241: out_data <= in_data241;
				'd242: out_data <= in_data242;
				'd243: out_data <= in_data243;
				'd244: out_data <= in_data244;
				'd245: out_data <= in_data245;
				'd246: out_data <= in_data246;
				'd247: out_data <= in_data247;
				'd248: out_data <= in_data248;
				'd249: out_data <= in_data249;
				'd250: out_data <= in_data250;
				'd251: out_data <= in_data251;
				'd252: out_data <= in_data252;
				'd253: out_data <= in_data253;
				'd254: out_data <= in_data254;
				'd255: out_data <= in_data255;
			endcase
		end
		else if (output_index==input_index && output_index!='d0) begin//finish dumping output
			out_data <= 'd0;
			out_valid <= 1'b0;
			dump_out_flag <= 1'b1;
		end
		else begin
			out_data <= 'd0;
			out_valid <= 1'b0;
		end
	end
	else begin
		out_data <= 'd0;
		out_valid <= 1'b0;
	end
end



/*
 * Combinational Block for exchaging elements of Bubble Sort
 */

reg			[7:0] temp_even1;
reg			[7:0] temp_even2;
reg			[7:0] temp_even3;
reg			[7:0] temp_even4;
reg			[7:0] temp_even5;
reg			[7:0] temp_even6;
reg			[7:0] temp_even7;
reg			[7:0] temp_even8;
reg			[7:0] temp_even9;
reg			[7:0] temp_even10;
reg			[7:0] temp_even11;
reg			[7:0] temp_even12;
reg			[7:0] temp_even13;
reg			[7:0] temp_even14;
reg			[7:0] temp_even15;
reg			[7:0] temp_even16;
reg			[7:0] temp_even17;
reg			[7:0] temp_even18;
reg			[7:0] temp_even19;
reg			[7:0] temp_even20;
reg			[7:0] temp_even21;
reg			[7:0] temp_even22;
reg			[7:0] temp_even23;
reg			[7:0] temp_even24;
reg			[7:0] temp_even25;
reg			[7:0] temp_even26;
reg			[7:0] temp_even27;
reg			[7:0] temp_even28;
reg			[7:0] temp_even29;
reg			[7:0] temp_even30;
reg			[7:0] temp_even31;
reg			[7:0] temp_even32;
reg			[7:0] temp_even33;
reg			[7:0] temp_even34;
reg			[7:0] temp_even35;
reg			[7:0] temp_even36;
reg			[7:0] temp_even37;
reg			[7:0] temp_even38;
reg			[7:0] temp_even39;
reg			[7:0] temp_even40;
reg			[7:0] temp_even41;
reg			[7:0] temp_even42;
reg			[7:0] temp_even43;
reg			[7:0] temp_even44;
reg			[7:0] temp_even45;
reg			[7:0] temp_even46;
reg			[7:0] temp_even47;
reg			[7:0] temp_even48;
reg			[7:0] temp_even49;
reg			[7:0] temp_even50;
reg			[7:0] temp_even51;
reg			[7:0] temp_even52;
reg			[7:0] temp_even53;
reg			[7:0] temp_even54;
reg			[7:0] temp_even55;
reg			[7:0] temp_even56;
reg			[7:0] temp_even57;
reg			[7:0] temp_even58;
reg			[7:0] temp_even59;
reg			[7:0] temp_even60;
reg			[7:0] temp_even61;
reg			[7:0] temp_even62;
reg			[7:0] temp_even63;
reg			[7:0] temp_even64;
reg			[7:0] temp_even65;
reg			[7:0] temp_even66;
reg			[7:0] temp_even67;
reg			[7:0] temp_even68;
reg			[7:0] temp_even69;
reg			[7:0] temp_even70;
reg			[7:0] temp_even71;
reg			[7:0] temp_even72;
reg			[7:0] temp_even73;
reg			[7:0] temp_even74;
reg			[7:0] temp_even75;
reg			[7:0] temp_even76;
reg			[7:0] temp_even77;
reg			[7:0] temp_even78;
reg			[7:0] temp_even79;
reg			[7:0] temp_even80;
reg			[7:0] temp_even81;
reg			[7:0] temp_even82;
reg			[7:0] temp_even83;
reg			[7:0] temp_even84;
reg			[7:0] temp_even85;
reg			[7:0] temp_even86;
reg			[7:0] temp_even87;
reg			[7:0] temp_even88;
reg			[7:0] temp_even89;
reg			[7:0] temp_even90;
reg			[7:0] temp_even91;
reg			[7:0] temp_even92;
reg			[7:0] temp_even93;
reg			[7:0] temp_even94;
reg			[7:0] temp_even95;
reg			[7:0] temp_even96;
reg			[7:0] temp_even97;
reg			[7:0] temp_even98;
reg			[7:0] temp_even99;
reg			[7:0] temp_even100;
reg			[7:0] temp_even101;
reg			[7:0] temp_even102;
reg			[7:0] temp_even103;
reg			[7:0] temp_even104;
reg			[7:0] temp_even105;
reg			[7:0] temp_even106;
reg			[7:0] temp_even107;
reg			[7:0] temp_even108;
reg			[7:0] temp_even109;
reg			[7:0] temp_even110;
reg			[7:0] temp_even111;
reg			[7:0] temp_even112;
reg			[7:0] temp_even113;
reg			[7:0] temp_even114;
reg			[7:0] temp_even115;
reg			[7:0] temp_even116;
reg			[7:0] temp_even117;
reg			[7:0] temp_even118;
reg			[7:0] temp_even119;
reg			[7:0] temp_even120;
reg			[7:0] temp_even121;
reg			[7:0] temp_even122;
reg			[7:0] temp_even123;
reg			[7:0] temp_even124;
reg			[7:0] temp_even125;
reg			[7:0] temp_even126;
reg			[7:0] temp_even127;
reg			[7:0] temp_even128;



reg			[7:0] temp_odd1;
reg			[7:0] temp_odd2;
reg			[7:0] temp_odd3;
reg			[7:0] temp_odd4;
reg			[7:0] temp_odd5;
reg			[7:0] temp_odd6;
reg			[7:0] temp_odd7;
reg			[7:0] temp_odd8;
reg			[7:0] temp_odd9;
reg			[7:0] temp_odd10;
reg			[7:0] temp_odd11;
reg			[7:0] temp_odd12;
reg			[7:0] temp_odd13;
reg			[7:0] temp_odd14;
reg			[7:0] temp_odd15;
reg			[7:0] temp_odd16;
reg			[7:0] temp_odd17;
reg			[7:0] temp_odd18;
reg			[7:0] temp_odd19;
reg			[7:0] temp_odd20;
reg			[7:0] temp_odd21;
reg			[7:0] temp_odd22;
reg			[7:0] temp_odd23;
reg			[7:0] temp_odd24;
reg			[7:0] temp_odd25;
reg			[7:0] temp_odd26;
reg			[7:0] temp_odd27;
reg			[7:0] temp_odd28;
reg			[7:0] temp_odd29;
reg			[7:0] temp_odd30;
reg			[7:0] temp_odd31;
reg			[7:0] temp_odd32;
reg			[7:0] temp_odd33;
reg			[7:0] temp_odd34;
reg			[7:0] temp_odd35;
reg			[7:0] temp_odd36;
reg			[7:0] temp_odd37;
reg			[7:0] temp_odd38;
reg			[7:0] temp_odd39;
reg			[7:0] temp_odd40;
reg			[7:0] temp_odd41;
reg			[7:0] temp_odd42;
reg			[7:0] temp_odd43;
reg			[7:0] temp_odd44;
reg			[7:0] temp_odd45;
reg			[7:0] temp_odd46;
reg			[7:0] temp_odd47;
reg			[7:0] temp_odd48;
reg			[7:0] temp_odd49;
reg			[7:0] temp_odd50;
reg			[7:0] temp_odd51;
reg			[7:0] temp_odd52;
reg			[7:0] temp_odd53;
reg			[7:0] temp_odd54;
reg			[7:0] temp_odd55;
reg			[7:0] temp_odd56;
reg			[7:0] temp_odd57;
reg			[7:0] temp_odd58;
reg			[7:0] temp_odd59;
reg			[7:0] temp_odd60;
reg			[7:0] temp_odd61;
reg			[7:0] temp_odd62;
reg			[7:0] temp_odd63;
reg			[7:0] temp_odd64;
reg			[7:0] temp_odd65;
reg			[7:0] temp_odd66;
reg			[7:0] temp_odd67;
reg			[7:0] temp_odd68;
reg			[7:0] temp_odd69;
reg			[7:0] temp_odd70;
reg			[7:0] temp_odd71;
reg			[7:0] temp_odd72;
reg			[7:0] temp_odd73;
reg			[7:0] temp_odd74;
reg			[7:0] temp_odd75;
reg			[7:0] temp_odd76;
reg			[7:0] temp_odd77;
reg			[7:0] temp_odd78;
reg			[7:0] temp_odd79;
reg			[7:0] temp_odd80;
reg			[7:0] temp_odd81;
reg			[7:0] temp_odd82;
reg			[7:0] temp_odd83;
reg			[7:0] temp_odd84;
reg			[7:0] temp_odd85;
reg			[7:0] temp_odd86;
reg			[7:0] temp_odd87;
reg			[7:0] temp_odd88;
reg			[7:0] temp_odd89;
reg			[7:0] temp_odd90;
reg			[7:0] temp_odd91;
reg			[7:0] temp_odd92;
reg			[7:0] temp_odd93;
reg			[7:0] temp_odd94;
reg			[7:0] temp_odd95;
reg			[7:0] temp_odd96;
reg			[7:0] temp_odd97;
reg			[7:0] temp_odd98;
reg			[7:0] temp_odd99;
reg			[7:0] temp_odd100;
reg			[7:0] temp_odd101;
reg			[7:0] temp_odd102;
reg			[7:0] temp_odd103;
reg			[7:0] temp_odd104;
reg			[7:0] temp_odd105;
reg			[7:0] temp_odd106;
reg			[7:0] temp_odd107;
reg			[7:0] temp_odd108;
reg			[7:0] temp_odd109;
reg			[7:0] temp_odd110;
reg			[7:0] temp_odd111;
reg			[7:0] temp_odd112;
reg			[7:0] temp_odd113;
reg			[7:0] temp_odd114;
reg			[7:0] temp_odd115;
reg			[7:0] temp_odd116;
reg			[7:0] temp_odd117;
reg			[7:0] temp_odd118;
reg			[7:0] temp_odd119;
reg			[7:0] temp_odd120;
reg			[7:0] temp_odd121;
reg			[7:0] temp_odd122;
reg			[7:0] temp_odd123;
reg			[7:0] temp_odd124;
reg			[7:0] temp_odd125;
reg			[7:0] temp_odd126;
reg			[7:0] temp_odd127;



always @(*) begin
	if (bubble_start_flag) begin
		if(outer_loop[0:0] == 1'b1) begin //odd
			if(in_data1 < in_data2) begin
				temp_odd1 = in_data1;
				in_data1 = in_data2;
				in_data2 = temp_odd1;
			end
			else begin
				temp_odd1 = 'd0;
			end
			if(in_data3 < in_data4) begin
				temp_odd2 = in_data3;
				in_data3 = in_data4;
				in_data4 = temp_odd2;
			end
			else begin
				temp_odd2 = 'd0;
			end
			if(in_data5 < in_data6) begin
				temp_odd3 = in_data5;
				in_data5 = in_data6;
				in_data6 = temp_odd3;
			end
			else begin
				temp_odd3 = 'd0;
			end
			if(in_data7 < in_data8) begin
				temp_odd4 = in_data7;
				in_data7 = in_data8;
				in_data8 = temp_odd4;
			end
			else begin
				temp_odd4 = 'd0;
			end
			if(in_data9 < in_data10) begin
				temp_odd5 = in_data9;
				in_data9 = in_data10;
				in_data10 = temp_odd5;
			end
			else begin
				temp_odd5 = 'd0;
			end
			if(in_data11 < in_data12) begin
				temp_odd6 = in_data11;
				in_data11 = in_data12;
				in_data12 = temp_odd6;
			end
			else begin
				temp_odd6 = 'd0;
			end
			if(in_data13 < in_data14) begin
				temp_odd7 = in_data13;
				in_data13 = in_data14;
				in_data14 = temp_odd7;
			end
			else begin
				temp_odd7 = 'd0;
			end
			if(in_data15 < in_data16) begin
				temp_odd8 = in_data15;
				in_data15 = in_data16;
				in_data16 = temp_odd8;
			end
			else begin
				temp_odd8 = 'd0;
			end
			if(in_data17 < in_data18) begin
				temp_odd9 = in_data17;
				in_data17 = in_data18;
				in_data18 = temp_odd9;
			end
			else begin
				temp_odd9 = 'd0;
			end
			if(in_data19 < in_data20) begin
				temp_odd10 = in_data19;
				in_data19 = in_data20;
				in_data20 = temp_odd10;
			end
			else begin
				temp_odd10 = 'd0;
			end
			if(in_data21 < in_data22) begin
				temp_odd11 = in_data21;
				in_data21 = in_data22;
				in_data22 = temp_odd11;
			end
			else begin
				temp_odd11 = 'd0;
			end
			if(in_data23 < in_data24) begin
				temp_odd12 = in_data23;
				in_data23 = in_data24;
				in_data24 = temp_odd12;
			end
			else begin
				temp_odd12 = 'd0;
			end
			if(in_data25 < in_data26) begin
				temp_odd13 = in_data25;
				in_data25 = in_data26;
				in_data26 = temp_odd13;
			end
			else begin
				temp_odd13 = 'd0;
			end
			if(in_data27 < in_data28) begin
				temp_odd14 = in_data27;
				in_data27 = in_data28;
				in_data28 = temp_odd14;
			end
			else begin
				temp_odd14 = 'd0;
			end
			if(in_data29 < in_data30) begin
				temp_odd15 = in_data29;
				in_data29 = in_data30;
				in_data30 = temp_odd15;
			end
			else begin
				temp_odd15 = 'd0;
			end
			if(in_data31 < in_data32) begin
				temp_odd16 = in_data31;
				in_data31 = in_data32;
				in_data32 = temp_odd16;
			end
			else begin
				temp_odd16 = 'd0;
			end
			if(in_data33 < in_data34) begin
				temp_odd17 = in_data33;
				in_data33 = in_data34;
				in_data34 = temp_odd17;
			end
			else begin
				temp_odd17 = 'd0;
			end
			if(in_data35 < in_data36) begin
				temp_odd18 = in_data35;
				in_data35 = in_data36;
				in_data36 = temp_odd18;
			end
			else begin
				temp_odd18 = 'd0;
			end
			if(in_data37 < in_data38) begin
				temp_odd19 = in_data37;
				in_data37 = in_data38;
				in_data38 = temp_odd19;
			end
			else begin
				temp_odd19 = 'd0;
			end
			if(in_data39 < in_data40) begin
				temp_odd20 = in_data39;
				in_data39 = in_data40;
				in_data40 = temp_odd20;
			end
			else begin
				temp_odd20 = 'd0;
			end
			if(in_data41 < in_data42) begin
				temp_odd21 = in_data41;
				in_data41 = in_data42;
				in_data42 = temp_odd21;
			end
			else begin
				temp_odd21 = 'd0;
			end
			if(in_data43 < in_data44) begin
				temp_odd22 = in_data43;
				in_data43 = in_data44;
				in_data44 = temp_odd22;
			end
			else begin
				temp_odd22 = 'd0;
			end
			if(in_data45 < in_data46) begin
				temp_odd23 = in_data45;
				in_data45 = in_data46;
				in_data46 = temp_odd23;
			end
			else begin
				temp_odd23 = 'd0;
			end
			if(in_data47 < in_data48) begin
				temp_odd24 = in_data47;
				in_data47 = in_data48;
				in_data48 = temp_odd24;
			end
			else begin
				temp_odd24 = 'd0;
			end
			if(in_data49 < in_data50) begin
				temp_odd25 = in_data49;
				in_data49 = in_data50;
				in_data50 = temp_odd25;
			end
			else begin
				temp_odd25 = 'd0;
			end
			if(in_data51 < in_data52) begin
				temp_odd26 = in_data51;
				in_data51 = in_data52;
				in_data52 = temp_odd26;
			end
			else begin
				temp_odd26 = 'd0;
			end
			if(in_data53 < in_data54) begin
				temp_odd27 = in_data53;
				in_data53 = in_data54;
				in_data54 = temp_odd27;
			end
			else begin
				temp_odd27 = 'd0;
			end
			if(in_data55 < in_data56) begin
				temp_odd28 = in_data55;
				in_data55 = in_data56;
				in_data56 = temp_odd28;
			end
			else begin
				temp_odd28 = 'd0;
			end
			if(in_data57 < in_data58) begin
				temp_odd29 = in_data57;
				in_data57 = in_data58;
				in_data58 = temp_odd29;
			end
			else begin
				temp_odd29 = 'd0;
			end
			if(in_data59 < in_data60) begin
				temp_odd30 = in_data59;
				in_data59 = in_data60;
				in_data60 = temp_odd30;
			end
			else begin
				temp_odd30 = 'd0;
			end
			if(in_data61 < in_data62) begin
				temp_odd31 = in_data61;
				in_data61 = in_data62;
				in_data62 = temp_odd31;
			end
			else begin
				temp_odd31 = 'd0;
			end
			if(in_data63 < in_data64) begin
				temp_odd32 = in_data63;
				in_data63 = in_data64;
				in_data64 = temp_odd32;
			end
			else begin
				temp_odd32 = 'd0;
			end
			if(in_data65 < in_data66) begin
				temp_odd33 = in_data65;
				in_data65 = in_data66;
				in_data66 = temp_odd33;
			end
			else begin
				temp_odd33 = 'd0;
			end
			if(in_data67 < in_data68) begin
				temp_odd34 = in_data67;
				in_data67 = in_data68;
				in_data68 = temp_odd34;
			end
			else begin
				temp_odd34 = 'd0;
			end
			if(in_data69 < in_data70) begin
				temp_odd35 = in_data69;
				in_data69 = in_data70;
				in_data70 = temp_odd35;
			end
			else begin
				temp_odd35 = 'd0;
			end
			if(in_data71 < in_data72) begin
				temp_odd36 = in_data71;
				in_data71 = in_data72;
				in_data72 = temp_odd36;
			end
			else begin
				temp_odd36 = 'd0;
			end
			if(in_data73 < in_data74) begin
				temp_odd37 = in_data73;
				in_data73 = in_data74;
				in_data74 = temp_odd37;
			end
			else begin
				temp_odd37 = 'd0;
			end
			if(in_data75 < in_data76) begin
				temp_odd38 = in_data75;
				in_data75 = in_data76;
				in_data76 = temp_odd38;
			end
			else begin
				temp_odd38 = 'd0;
			end
			if(in_data77 < in_data78) begin
				temp_odd39 = in_data77;
				in_data77 = in_data78;
				in_data78 = temp_odd39;
			end
			else begin
				temp_odd39 = 'd0;
			end
			if(in_data79 < in_data80) begin
				temp_odd40 = in_data79;
				in_data79 = in_data80;
				in_data80 = temp_odd40;
			end
			else begin
				temp_odd40 = 'd0;
			end
			if(in_data81 < in_data82) begin
				temp_odd41 = in_data81;
				in_data81 = in_data82;
				in_data82 = temp_odd41;
			end
			else begin
				temp_odd41 = 'd0;
			end
			if(in_data83 < in_data84) begin
				temp_odd42 = in_data83;
				in_data83 = in_data84;
				in_data84 = temp_odd42;
			end
			else begin
				temp_odd42 = 'd0;
			end
			if(in_data85 < in_data86) begin
				temp_odd43 = in_data85;
				in_data85 = in_data86;
				in_data86 = temp_odd43;
			end
			else begin
				temp_odd43 = 'd0;
			end
			if(in_data87 < in_data88) begin
				temp_odd44 = in_data87;
				in_data87 = in_data88;
				in_data88 = temp_odd44;
			end
			else begin
				temp_odd44 = 'd0;
			end
			if(in_data89 < in_data90) begin
				temp_odd45 = in_data89;
				in_data89 = in_data90;
				in_data90 = temp_odd45;
			end
			else begin
				temp_odd45 = 'd0;
			end
			if(in_data91 < in_data92) begin
				temp_odd46 = in_data91;
				in_data91 = in_data92;
				in_data92 = temp_odd46;
			end
			else begin
				temp_odd46 = 'd0;
			end
			if(in_data93 < in_data94) begin
				temp_odd47 = in_data93;
				in_data93 = in_data94;
				in_data94 = temp_odd47;
			end
			else begin
				temp_odd47 = 'd0;
			end
			if(in_data95 < in_data96) begin
				temp_odd48 = in_data95;
				in_data95 = in_data96;
				in_data96 = temp_odd48;
			end
			else begin
				temp_odd48 = 'd0;
			end
			if(in_data97 < in_data98) begin
				temp_odd49 = in_data97;
				in_data97 = in_data98;
				in_data98 = temp_odd49;
			end
			else begin
				temp_odd49 = 'd0;
			end
			if(in_data99 < in_data100) begin
				temp_odd50 = in_data99;
				in_data99 = in_data100;
				in_data100 = temp_odd50;
			end
			else begin
				temp_odd50 = 'd0;
			end
			if(in_data101 < in_data102) begin
				temp_odd51 = in_data101;
				in_data101 = in_data102;
				in_data102 = temp_odd51;
			end
			else begin
				temp_odd51 = 'd0;
			end
			if(in_data103 < in_data104) begin
				temp_odd52 = in_data103;
				in_data103 = in_data104;
				in_data104 = temp_odd52;
			end
			else begin
				temp_odd52 = 'd0;
			end
			if(in_data105 < in_data106) begin
				temp_odd53 = in_data105;
				in_data105 = in_data106;
				in_data106 = temp_odd53;
			end
			else begin
				temp_odd53 = 'd0;
			end
			if(in_data107 < in_data108) begin
				temp_odd54 = in_data107;
				in_data107 = in_data108;
				in_data108 = temp_odd54;
			end
			else begin
				temp_odd54 = 'd0;
			end
			if(in_data109 < in_data110) begin
				temp_odd55 = in_data109;
				in_data109 = in_data110;
				in_data110 = temp_odd55;
			end
			else begin
				temp_odd55 = 'd0;
			end
			if(in_data111 < in_data112) begin
				temp_odd56 = in_data111;
				in_data111 = in_data112;
				in_data112 = temp_odd56;
			end
			else begin
				temp_odd56 = 'd0;
			end
			if(in_data113 < in_data114) begin
				temp_odd57 = in_data113;
				in_data113 = in_data114;
				in_data114 = temp_odd57;
			end
			else begin
				temp_odd57 = 'd0;
			end
			if(in_data115 < in_data116) begin
				temp_odd58 = in_data115;
				in_data115 = in_data116;
				in_data116 = temp_odd58;
			end
			else begin
				temp_odd58 = 'd0;
			end
			if(in_data117 < in_data118) begin
				temp_odd59 = in_data117;
				in_data117 = in_data118;
				in_data118 = temp_odd59;
			end
			else begin
				temp_odd59 = 'd0;
			end
			if(in_data119 < in_data120) begin
				temp_odd60 = in_data119;
				in_data119 = in_data120;
				in_data120 = temp_odd60;
			end
			else begin
				temp_odd60 = 'd0;
			end
			if(in_data121 < in_data122) begin
				temp_odd61 = in_data121;
				in_data121 = in_data122;
				in_data122 = temp_odd61;
			end
			else begin
				temp_odd61 = 'd0;
			end
			if(in_data123 < in_data124) begin
				temp_odd62 = in_data123;
				in_data123 = in_data124;
				in_data124 = temp_odd62;
			end
			else begin
				temp_odd62 = 'd0;
			end
			if(in_data125 < in_data126) begin
				temp_odd63 = in_data125;
				in_data125 = in_data126;
				in_data126 = temp_odd63;
			end
			else begin
				temp_odd63 = 'd0;
			end
			if(in_data127 < in_data128) begin
				temp_odd64 = in_data127;
				in_data127 = in_data128;
				in_data128 = temp_odd64;
			end
			else begin
				temp_odd64 = 'd0;
			end
			if(in_data129 < in_data130) begin
				temp_odd65 = in_data129;
				in_data129 = in_data130;
				in_data130 = temp_odd65;
			end
			else begin
				temp_odd65 = 'd0;
			end
			if(in_data131 < in_data132) begin
				temp_odd66 = in_data131;
				in_data131 = in_data132;
				in_data132 = temp_odd66;
			end
			else begin
				temp_odd66 = 'd0;
			end
			if(in_data133 < in_data134) begin
				temp_odd67 = in_data133;
				in_data133 = in_data134;
				in_data134 = temp_odd67;
			end
			else begin
				temp_odd67 = 'd0;
			end
			if(in_data135 < in_data136) begin
				temp_odd68 = in_data135;
				in_data135 = in_data136;
				in_data136 = temp_odd68;
			end
			else begin
				temp_odd68 = 'd0;
			end
			if(in_data137 < in_data138) begin
				temp_odd69 = in_data137;
				in_data137 = in_data138;
				in_data138 = temp_odd69;
			end
			else begin
				temp_odd69 = 'd0;
			end
			if(in_data139 < in_data140) begin
				temp_odd70 = in_data139;
				in_data139 = in_data140;
				in_data140 = temp_odd70;
			end
			else begin
				temp_odd70 = 'd0;
			end
			if(in_data141 < in_data142) begin
				temp_odd71 = in_data141;
				in_data141 = in_data142;
				in_data142 = temp_odd71;
			end
			else begin
				temp_odd71 = 'd0;
			end
			if(in_data143 < in_data144) begin
				temp_odd72 = in_data143;
				in_data143 = in_data144;
				in_data144 = temp_odd72;
			end
			else begin
				temp_odd72 = 'd0;
			end
			if(in_data145 < in_data146) begin
				temp_odd73 = in_data145;
				in_data145 = in_data146;
				in_data146 = temp_odd73;
			end
			else begin
				temp_odd73 = 'd0;
			end
			if(in_data147 < in_data148) begin
				temp_odd74 = in_data147;
				in_data147 = in_data148;
				in_data148 = temp_odd74;
			end
			else begin
				temp_odd74 = 'd0;
			end
			if(in_data149 < in_data150) begin
				temp_odd75 = in_data149;
				in_data149 = in_data150;
				in_data150 = temp_odd75;
			end
			else begin
				temp_odd75 = 'd0;
			end
			if(in_data151 < in_data152) begin
				temp_odd76 = in_data151;
				in_data151 = in_data152;
				in_data152 = temp_odd76;
			end
			else begin
				temp_odd76 = 'd0;
			end
			if(in_data153 < in_data154) begin
				temp_odd77 = in_data153;
				in_data153 = in_data154;
				in_data154 = temp_odd77;
			end
			else begin
				temp_odd77 = 'd0;
			end
			if(in_data155 < in_data156) begin
				temp_odd78 = in_data155;
				in_data155 = in_data156;
				in_data156 = temp_odd78;
			end
			else begin
				temp_odd78 = 'd0;
			end
			if(in_data157 < in_data158) begin
				temp_odd79 = in_data157;
				in_data157 = in_data158;
				in_data158 = temp_odd79;
			end
			else begin
				temp_odd79 = 'd0;
			end
			if(in_data159 < in_data160) begin
				temp_odd80 = in_data159;
				in_data159 = in_data160;
				in_data160 = temp_odd80;
			end
			else begin
				temp_odd80 = 'd0;
			end
			if(in_data161 < in_data162) begin
				temp_odd81 = in_data161;
				in_data161 = in_data162;
				in_data162 = temp_odd81;
			end
			else begin
				temp_odd81 = 'd0;
			end
			if(in_data163 < in_data164) begin
				temp_odd82 = in_data163;
				in_data163 = in_data164;
				in_data164 = temp_odd82;
			end
			else begin
				temp_odd82 = 'd0;
			end
			if(in_data165 < in_data166) begin
				temp_odd83 = in_data165;
				in_data165 = in_data166;
				in_data166 = temp_odd83;
			end
			else begin
				temp_odd83 = 'd0;
			end
			if(in_data167 < in_data168) begin
				temp_odd84 = in_data167;
				in_data167 = in_data168;
				in_data168 = temp_odd84;
			end
			else begin
				temp_odd84 = 'd0;
			end
			if(in_data169 < in_data170) begin
				temp_odd85 = in_data169;
				in_data169 = in_data170;
				in_data170 = temp_odd85;
			end
			else begin
				temp_odd85 = 'd0;
			end
			if(in_data171 < in_data172) begin
				temp_odd86 = in_data171;
				in_data171 = in_data172;
				in_data172 = temp_odd86;
			end
			else begin
				temp_odd86 = 'd0;
			end
			if(in_data173 < in_data174) begin
				temp_odd87 = in_data173;
				in_data173 = in_data174;
				in_data174 = temp_odd87;
			end
			else begin
				temp_odd87 = 'd0;
			end
			if(in_data175 < in_data176) begin
				temp_odd88 = in_data175;
				in_data175 = in_data176;
				in_data176 = temp_odd88;
			end
			else begin
				temp_odd88 = 'd0;
			end
			if(in_data177 < in_data178) begin
				temp_odd89 = in_data177;
				in_data177 = in_data178;
				in_data178 = temp_odd89;
			end
			else begin
				temp_odd89 = 'd0;
			end
			if(in_data179 < in_data180) begin
				temp_odd90 = in_data179;
				in_data179 = in_data180;
				in_data180 = temp_odd90;
			end
			else begin
				temp_odd90 = 'd0;
			end
			if(in_data181 < in_data182) begin
				temp_odd91 = in_data181;
				in_data181 = in_data182;
				in_data182 = temp_odd91;
			end
			else begin
				temp_odd91 = 'd0;
			end
			if(in_data183 < in_data184) begin
				temp_odd92 = in_data183;
				in_data183 = in_data184;
				in_data184 = temp_odd92;
			end
			else begin
				temp_odd92 = 'd0;
			end
			if(in_data185 < in_data186) begin
				temp_odd93 = in_data185;
				in_data185 = in_data186;
				in_data186 = temp_odd93;
			end
			else begin
				temp_odd93 = 'd0;
			end
			if(in_data187 < in_data188) begin
				temp_odd94 = in_data187;
				in_data187 = in_data188;
				in_data188 = temp_odd94;
			end
			else begin
				temp_odd94 = 'd0;
			end
			if(in_data189 < in_data190) begin
				temp_odd95 = in_data189;
				in_data189 = in_data190;
				in_data190 = temp_odd95;
			end
			else begin
				temp_odd95 = 'd0;
			end
			if(in_data191 < in_data192) begin
				temp_odd96 = in_data191;
				in_data191 = in_data192;
				in_data192 = temp_odd96;
			end
			else begin
				temp_odd96 = 'd0;
			end
			if(in_data193 < in_data194) begin
				temp_odd97 = in_data193;
				in_data193 = in_data194;
				in_data194 = temp_odd97;
			end
			else begin
				temp_odd97 = 'd0;
			end
			if(in_data195 < in_data196) begin
				temp_odd98 = in_data195;
				in_data195 = in_data196;
				in_data196 = temp_odd98;
			end
			else begin
				temp_odd98 = 'd0;
			end
			if(in_data197 < in_data198) begin
				temp_odd99 = in_data197;
				in_data197 = in_data198;
				in_data198 = temp_odd99;
			end
			else begin
				temp_odd99 = 'd0;
			end
			if(in_data199 < in_data200) begin
				temp_odd100 = in_data199;
				in_data199 = in_data200;
				in_data200 = temp_odd100;
			end
			else begin
				temp_odd100 = 'd0;
			end
			if(in_data201 < in_data202) begin
				temp_odd101 = in_data201;
				in_data201 = in_data202;
				in_data202 = temp_odd101;
			end
			else begin
				temp_odd101 = 'd0;
			end
			if(in_data203 < in_data204) begin
				temp_odd102 = in_data203;
				in_data203 = in_data204;
				in_data204 = temp_odd102;
			end
			else begin
				temp_odd102 = 'd0;
			end
			if(in_data205 < in_data206) begin
				temp_odd103 = in_data205;
				in_data205 = in_data206;
				in_data206 = temp_odd103;
			end
			else begin
				temp_odd103 = 'd0;
			end
			if(in_data207 < in_data208) begin
				temp_odd104 = in_data207;
				in_data207 = in_data208;
				in_data208 = temp_odd104;
			end
			else begin
				temp_odd104 = 'd0;
			end
			if(in_data209 < in_data210) begin
				temp_odd105 = in_data209;
				in_data209 = in_data210;
				in_data210 = temp_odd105;
			end
			else begin
				temp_odd105 = 'd0;
			end
			if(in_data211 < in_data212) begin
				temp_odd106 = in_data211;
				in_data211 = in_data212;
				in_data212 = temp_odd106;
			end
			else begin
				temp_odd106 = 'd0;
			end
			if(in_data213 < in_data214) begin
				temp_odd107 = in_data213;
				in_data213 = in_data214;
				in_data214 = temp_odd107;
			end
			else begin
				temp_odd107 = 'd0;
			end
			if(in_data215 < in_data216) begin
				temp_odd108 = in_data215;
				in_data215 = in_data216;
				in_data216 = temp_odd108;
			end
			else begin
				temp_odd108 = 'd0;
			end
			if(in_data217 < in_data218) begin
				temp_odd109 = in_data217;
				in_data217 = in_data218;
				in_data218 = temp_odd109;
			end
			else begin
				temp_odd109 = 'd0;
			end
			if(in_data219 < in_data220) begin
				temp_odd110 = in_data219;
				in_data219 = in_data220;
				in_data220 = temp_odd110;
			end
			else begin
				temp_odd110 = 'd0;
			end
			if(in_data221 < in_data222) begin
				temp_odd111 = in_data221;
				in_data221 = in_data222;
				in_data222 = temp_odd111;
			end
			else begin
				temp_odd111 = 'd0;
			end
			if(in_data223 < in_data224) begin
				temp_odd112 = in_data223;
				in_data223 = in_data224;
				in_data224 = temp_odd112;
			end
			else begin
				temp_odd112 = 'd0;
			end
			if(in_data225 < in_data226) begin
				temp_odd113 = in_data225;
				in_data225 = in_data226;
				in_data226 = temp_odd113;
			end
			else begin
				temp_odd113 = 'd0;
			end
			if(in_data227 < in_data228) begin
				temp_odd114 = in_data227;
				in_data227 = in_data228;
				in_data228 = temp_odd114;
			end
			else begin
				temp_odd114 = 'd0;
			end
			if(in_data229 < in_data230) begin
				temp_odd115 = in_data229;
				in_data229 = in_data230;
				in_data230 = temp_odd115;
			end
			else begin
				temp_odd115 = 'd0;
			end
			if(in_data231 < in_data232) begin
				temp_odd116 = in_data231;
				in_data231 = in_data232;
				in_data232 = temp_odd116;
			end
			else begin
				temp_odd116 = 'd0;
			end
			if(in_data233 < in_data234) begin
				temp_odd117 = in_data233;
				in_data233 = in_data234;
				in_data234 = temp_odd117;
			end
			else begin
				temp_odd117 = 'd0;
			end
			if(in_data235 < in_data236) begin
				temp_odd118 = in_data235;
				in_data235 = in_data236;
				in_data236 = temp_odd118;
			end
			else begin
				temp_odd118 = 'd0;
			end
			if(in_data237 < in_data238) begin
				temp_odd119 = in_data237;
				in_data237 = in_data238;
				in_data238 = temp_odd119;
			end
			else begin
				temp_odd119 = 'd0;
			end
			if(in_data239 < in_data240) begin
				temp_odd120 = in_data239;
				in_data239 = in_data240;
				in_data240 = temp_odd120;
			end
			else begin
				temp_odd120 = 'd0;
			end
			if(in_data241 < in_data242) begin
				temp_odd121 = in_data241;
				in_data241 = in_data242;
				in_data242 = temp_odd121;
			end
			else begin
				temp_odd121 = 'd0;
			end
			if(in_data243 < in_data244) begin
				temp_odd122 = in_data243;
				in_data243 = in_data244;
				in_data244 = temp_odd122;
			end
			else begin
				temp_odd122 = 'd0;
			end
			if(in_data245 < in_data246) begin
				temp_odd123 = in_data245;
				in_data245 = in_data246;
				in_data246 = temp_odd123;
			end
			else begin
				temp_odd123 = 'd0;
			end
			if(in_data247 < in_data248) begin
				temp_odd124 = in_data247;
				in_data247 = in_data248;
				in_data248 = temp_odd124;
			end
			else begin
				temp_odd124 = 'd0;
			end
			if(in_data249 < in_data250) begin
				temp_odd125 = in_data249;
				in_data249 = in_data250;
				in_data250 = temp_odd125;
			end
			else begin
				temp_odd125 = 'd0;
			end
			if(in_data251 < in_data252) begin
				temp_odd126 = in_data251;
				in_data251 = in_data252;
				in_data252 = temp_odd126;
			end
			else begin
				temp_odd126 = 'd0;
			end
			if(in_data253 < in_data254) begin
				temp_odd127 = in_data253;
				in_data253 = in_data254;
				in_data254 = temp_odd127;
			end
			else begin
				temp_odd127 = 'd0;
			end
		end
		else begin //even
			if (in_data0 < in_data1) begin
				temp_even1 = in_data0;
				in_data0 = in_data1;
				in_data1 = temp_even1;
			end
			else begin
				temp_even1 = 'd0;
			end
			if (in_data2 < in_data3) begin
				temp_even2 = in_data2;
				in_data2 = in_data3;
				in_data3 = temp_even2;
			end
			else begin
				temp_even2 = 'd0;
			end
			if (in_data4 < in_data5) begin
				temp_even3 = in_data4;
				in_data4 = in_data5;
				in_data5 = temp_even3;
			end
			else begin
				temp_even3 = 'd0;
			end
			if (in_data6 < in_data7) begin
				temp_even4 = in_data6;
				in_data6 = in_data7;
				in_data7 = temp_even4;
			end
			else begin
				temp_even4 = 'd0;
			end
			if (in_data8 < in_data9) begin
				temp_even5 = in_data8;
				in_data8 = in_data9;
				in_data9 = temp_even5;
			end
			else begin
				temp_even5 = 'd0;
			end
			if (in_data10 < in_data11) begin
				temp_even6 = in_data10;
				in_data10 = in_data11;
				in_data11 = temp_even6;
			end
			else begin
				temp_even6 = 'd0;
			end
			if (in_data12 < in_data13) begin
				temp_even7 = in_data12;
				in_data12 = in_data13;
				in_data13 = temp_even7;
			end
			else begin
				temp_even7 = 'd0;
			end
			if (in_data14 < in_data15) begin
				temp_even8 = in_data14;
				in_data14 = in_data15;
				in_data15 = temp_even8;
			end
			else begin
				temp_even8 = 'd0;
			end
			if (in_data16 < in_data17) begin
				temp_even9 = in_data16;
				in_data16 = in_data17;
				in_data17 = temp_even9;
			end
			else begin
				temp_even9 = 'd0;
			end
			if (in_data18 < in_data19) begin
				temp_even10 = in_data18;
				in_data18 = in_data19;
				in_data19 = temp_even10;
			end
			else begin
				temp_even10 = 'd0;
			end
			if (in_data20 < in_data21) begin
				temp_even11 = in_data20;
				in_data20 = in_data21;
				in_data21 = temp_even11;
			end
			else begin
				temp_even11 = 'd0;
			end
			if (in_data22 < in_data23) begin
				temp_even12 = in_data22;
				in_data22 = in_data23;
				in_data23 = temp_even12;
			end
			else begin
				temp_even12 = 'd0;
			end
			if (in_data24 < in_data25) begin
				temp_even13 = in_data24;
				in_data24 = in_data25;
				in_data25 = temp_even13;
			end
			else begin
				temp_even13 = 'd0;
			end
			if (in_data26 < in_data27) begin
				temp_even14 = in_data26;
				in_data26 = in_data27;
				in_data27 = temp_even14;
			end
			else begin
				temp_even14 = 'd0;
			end
			if (in_data28 < in_data29) begin
				temp_even15 = in_data28;
				in_data28 = in_data29;
				in_data29 = temp_even15;
			end
			else begin
				temp_even15 = 'd0;
			end
			if (in_data30 < in_data31) begin
				temp_even16 = in_data30;
				in_data30 = in_data31;
				in_data31 = temp_even16;
			end
			else begin
				temp_even16 = 'd0;
			end
			if (in_data32 < in_data33) begin
				temp_even17 = in_data32;
				in_data32 = in_data33;
				in_data33 = temp_even17;
			end
			else begin
				temp_even17 = 'd0;
			end
			if (in_data34 < in_data35) begin
				temp_even18 = in_data34;
				in_data34 = in_data35;
				in_data35 = temp_even18;
			end
			else begin
				temp_even18 = 'd0;
			end
			if (in_data36 < in_data37) begin
				temp_even19 = in_data36;
				in_data36 = in_data37;
				in_data37 = temp_even19;
			end
			else begin
				temp_even19 = 'd0;
			end
			if (in_data38 < in_data39) begin
				temp_even20 = in_data38;
				in_data38 = in_data39;
				in_data39 = temp_even20;
			end
			else begin
				temp_even20 = 'd0;
			end
			if (in_data40 < in_data41) begin
				temp_even21 = in_data40;
				in_data40 = in_data41;
				in_data41 = temp_even21;
			end
			else begin
				temp_even21 = 'd0;
			end
			if (in_data42 < in_data43) begin
				temp_even22 = in_data42;
				in_data42 = in_data43;
				in_data43 = temp_even22;
			end
			else begin
				temp_even22 = 'd0;
			end
			if (in_data44 < in_data45) begin
				temp_even23 = in_data44;
				in_data44 = in_data45;
				in_data45 = temp_even23;
			end
			else begin
				temp_even23 = 'd0;
			end
			if (in_data46 < in_data47) begin
				temp_even24 = in_data46;
				in_data46 = in_data47;
				in_data47 = temp_even24;
			end
			else begin
				temp_even24 = 'd0;
			end
			if (in_data48 < in_data49) begin
				temp_even25 = in_data48;
				in_data48 = in_data49;
				in_data49 = temp_even25;
			end
			else begin
				temp_even25 = 'd0;
			end
			if (in_data50 < in_data51) begin
				temp_even26 = in_data50;
				in_data50 = in_data51;
				in_data51 = temp_even26;
			end
			else begin
				temp_even26 = 'd0;
			end
			if (in_data52 < in_data53) begin
				temp_even27 = in_data52;
				in_data52 = in_data53;
				in_data53 = temp_even27;
			end
			else begin
				temp_even27 = 'd0;
			end
			if (in_data54 < in_data55) begin
				temp_even28 = in_data54;
				in_data54 = in_data55;
				in_data55 = temp_even28;
			end
			else begin
				temp_even28 = 'd0;
			end
			if (in_data56 < in_data57) begin
				temp_even29 = in_data56;
				in_data56 = in_data57;
				in_data57 = temp_even29;
			end
			else begin
				temp_even29 = 'd0;
			end
			if (in_data58 < in_data59) begin
				temp_even30 = in_data58;
				in_data58 = in_data59;
				in_data59 = temp_even30;
			end
			else begin
				temp_even30 = 'd0;
			end
			if (in_data60 < in_data61) begin
				temp_even31 = in_data60;
				in_data60 = in_data61;
				in_data61 = temp_even31;
			end
			else begin
				temp_even31 = 'd0;
			end
			if (in_data62 < in_data63) begin
				temp_even32 = in_data62;
				in_data62 = in_data63;
				in_data63 = temp_even32;
			end
			else begin
				temp_even32 = 'd0;
			end
			if (in_data64 < in_data65) begin
				temp_even33 = in_data64;
				in_data64 = in_data65;
				in_data65 = temp_even33;
			end
			else begin
				temp_even33 = 'd0;
			end
			if (in_data66 < in_data67) begin
				temp_even34 = in_data66;
				in_data66 = in_data67;
				in_data67 = temp_even34;
			end
			else begin
				temp_even34 = 'd0;
			end
			if (in_data68 < in_data69) begin
				temp_even35 = in_data68;
				in_data68 = in_data69;
				in_data69 = temp_even35;
			end
			else begin
				temp_even35 = 'd0;
			end
			if (in_data70 < in_data71) begin
				temp_even36 = in_data70;
				in_data70 = in_data71;
				in_data71 = temp_even36;
			end
			else begin
				temp_even36 = 'd0;
			end
			if (in_data72 < in_data73) begin
				temp_even37 = in_data72;
				in_data72 = in_data73;
				in_data73 = temp_even37;
			end
			else begin
				temp_even37 = 'd0;
			end
			if (in_data74 < in_data75) begin
				temp_even38 = in_data74;
				in_data74 = in_data75;
				in_data75 = temp_even38;
			end
			else begin
				temp_even38 = 'd0;
			end
			if (in_data76 < in_data77) begin
				temp_even39 = in_data76;
				in_data76 = in_data77;
				in_data77 = temp_even39;
			end
			else begin
				temp_even39 = 'd0;
			end
			if (in_data78 < in_data79) begin
				temp_even40 = in_data78;
				in_data78 = in_data79;
				in_data79 = temp_even40;
			end
			else begin
				temp_even40 = 'd0;
			end
			if (in_data80 < in_data81) begin
				temp_even41 = in_data80;
				in_data80 = in_data81;
				in_data81 = temp_even41;
			end
			else begin
				temp_even41 = 'd0;
			end
			if (in_data82 < in_data83) begin
				temp_even42 = in_data82;
				in_data82 = in_data83;
				in_data83 = temp_even42;
			end
			else begin
				temp_even42 = 'd0;
			end
			if (in_data84 < in_data85) begin
				temp_even43 = in_data84;
				in_data84 = in_data85;
				in_data85 = temp_even43;
			end
			else begin
				temp_even43 = 'd0;
			end
			if (in_data86 < in_data87) begin
				temp_even44 = in_data86;
				in_data86 = in_data87;
				in_data87 = temp_even44;
			end
			else begin
				temp_even44 = 'd0;
			end
			if (in_data88 < in_data89) begin
				temp_even45 = in_data88;
				in_data88 = in_data89;
				in_data89 = temp_even45;
			end
			else begin
				temp_even45 = 'd0;
			end
			if (in_data90 < in_data91) begin
				temp_even46 = in_data90;
				in_data90 = in_data91;
				in_data91 = temp_even46;
			end
			else begin
				temp_even46 = 'd0;
			end
			if (in_data92 < in_data93) begin
				temp_even47 = in_data92;
				in_data92 = in_data93;
				in_data93 = temp_even47;
			end
			else begin
				temp_even47 = 'd0;
			end
			if (in_data94 < in_data95) begin
				temp_even48 = in_data94;
				in_data94 = in_data95;
				in_data95 = temp_even48;
			end
			else begin
				temp_even48 = 'd0;
			end
			if (in_data96 < in_data97) begin
				temp_even49 = in_data96;
				in_data96 = in_data97;
				in_data97 = temp_even49;
			end
			else begin
				temp_even49 = 'd0;
			end
			if (in_data98 < in_data99) begin
				temp_even50 = in_data98;
				in_data98 = in_data99;
				in_data99 = temp_even50;
			end
			else begin
				temp_even50 = 'd0;
			end
			if (in_data100 < in_data101) begin
				temp_even51 = in_data100;
				in_data100 = in_data101;
				in_data101 = temp_even51;
			end
			else begin
				temp_even51 = 'd0;
			end
			if (in_data102 < in_data103) begin
				temp_even52 = in_data102;
				in_data102 = in_data103;
				in_data103 = temp_even52;
			end
			else begin
				temp_even52 = 'd0;
			end
			if (in_data104 < in_data105) begin
				temp_even53 = in_data104;
				in_data104 = in_data105;
				in_data105 = temp_even53;
			end
			else begin
				temp_even53 = 'd0;
			end
			if (in_data106 < in_data107) begin
				temp_even54 = in_data106;
				in_data106 = in_data107;
				in_data107 = temp_even54;
			end
			else begin
				temp_even54 = 'd0;
			end
			if (in_data108 < in_data109) begin
				temp_even55 = in_data108;
				in_data108 = in_data109;
				in_data109 = temp_even55;
			end
			else begin
				temp_even55 = 'd0;
			end
			if (in_data110 < in_data111) begin
				temp_even56 = in_data110;
				in_data110 = in_data111;
				in_data111 = temp_even56;
			end
			else begin
				temp_even56 = 'd0;
			end
			if (in_data112 < in_data113) begin
				temp_even57 = in_data112;
				in_data112 = in_data113;
				in_data113 = temp_even57;
			end
			else begin
				temp_even57 = 'd0;
			end
			if (in_data114 < in_data115) begin
				temp_even58 = in_data114;
				in_data114 = in_data115;
				in_data115 = temp_even58;
			end
			else begin
				temp_even58 = 'd0;
			end
			if (in_data116 < in_data117) begin
				temp_even59 = in_data116;
				in_data116 = in_data117;
				in_data117 = temp_even59;
			end
			else begin
				temp_even59 = 'd0;
			end
			if (in_data118 < in_data119) begin
				temp_even60 = in_data118;
				in_data118 = in_data119;
				in_data119 = temp_even60;
			end
			else begin
				temp_even60 = 'd0;
			end
			if (in_data120 < in_data121) begin
				temp_even61 = in_data120;
				in_data120 = in_data121;
				in_data121 = temp_even61;
			end
			else begin
				temp_even61 = 'd0;
			end
			if (in_data122 < in_data123) begin
				temp_even62 = in_data122;
				in_data122 = in_data123;
				in_data123 = temp_even62;
			end
			else begin
				temp_even62 = 'd0;
			end
			if (in_data124 < in_data125) begin
				temp_even63 = in_data124;
				in_data124 = in_data125;
				in_data125 = temp_even63;
			end
			else begin
				temp_even63 = 'd0;
			end
			if (in_data126 < in_data127) begin
				temp_even64 = in_data126;
				in_data126 = in_data127;
				in_data127 = temp_even64;
			end
			else begin
				temp_even64 = 'd0;
			end
			if (in_data128 < in_data129) begin
				temp_even65 = in_data128;
				in_data128 = in_data129;
				in_data129 = temp_even65;
			end
			else begin
				temp_even65 = 'd0;
			end
			if (in_data130 < in_data131) begin
				temp_even66 = in_data130;
				in_data130 = in_data131;
				in_data131 = temp_even66;
			end
			else begin
				temp_even66 = 'd0;
			end
			if (in_data132 < in_data133) begin
				temp_even67 = in_data132;
				in_data132 = in_data133;
				in_data133 = temp_even67;
			end
			else begin
				temp_even67 = 'd0;
			end
			if (in_data134 < in_data135) begin
				temp_even68 = in_data134;
				in_data134 = in_data135;
				in_data135 = temp_even68;
			end
			else begin
				temp_even68 = 'd0;
			end
			if (in_data136 < in_data137) begin
				temp_even69 = in_data136;
				in_data136 = in_data137;
				in_data137 = temp_even69;
			end
			else begin
				temp_even69 = 'd0;
			end
			if (in_data138 < in_data139) begin
				temp_even70 = in_data138;
				in_data138 = in_data139;
				in_data139 = temp_even70;
			end
			else begin
				temp_even70 = 'd0;
			end
			if (in_data140 < in_data141) begin
				temp_even71 = in_data140;
				in_data140 = in_data141;
				in_data141 = temp_even71;
			end
			else begin
				temp_even71 = 'd0;
			end
			if (in_data142 < in_data143) begin
				temp_even72 = in_data142;
				in_data142 = in_data143;
				in_data143 = temp_even72;
			end
			else begin
				temp_even72 = 'd0;
			end
			if (in_data144 < in_data145) begin
				temp_even73 = in_data144;
				in_data144 = in_data145;
				in_data145 = temp_even73;
			end
			else begin
				temp_even73 = 'd0;
			end
			if (in_data146 < in_data147) begin
				temp_even74 = in_data146;
				in_data146 = in_data147;
				in_data147 = temp_even74;
			end
			else begin
				temp_even74 = 'd0;
			end
			if (in_data148 < in_data149) begin
				temp_even75 = in_data148;
				in_data148 = in_data149;
				in_data149 = temp_even75;
			end
			else begin
				temp_even75 = 'd0;
			end
			if (in_data150 < in_data151) begin
				temp_even76 = in_data150;
				in_data150 = in_data151;
				in_data151 = temp_even76;
			end
			else begin
				temp_even76 = 'd0;
			end
			if (in_data152 < in_data153) begin
				temp_even77 = in_data152;
				in_data152 = in_data153;
				in_data153 = temp_even77;
			end
			else begin
				temp_even77 = 'd0;
			end
			if (in_data154 < in_data155) begin
				temp_even78 = in_data154;
				in_data154 = in_data155;
				in_data155 = temp_even78;
			end
			else begin
				temp_even78 = 'd0;
			end
			if (in_data156 < in_data157) begin
				temp_even79 = in_data156;
				in_data156 = in_data157;
				in_data157 = temp_even79;
			end
			else begin
				temp_even79 = 'd0;
			end
			if (in_data158 < in_data159) begin
				temp_even80 = in_data158;
				in_data158 = in_data159;
				in_data159 = temp_even80;
			end
			else begin
				temp_even80 = 'd0;
			end
			if (in_data160 < in_data161) begin
				temp_even81 = in_data160;
				in_data160 = in_data161;
				in_data161 = temp_even81;
			end
			else begin
				temp_even81 = 'd0;
			end
			if (in_data162 < in_data163) begin
				temp_even82 = in_data162;
				in_data162 = in_data163;
				in_data163 = temp_even82;
			end
			else begin
				temp_even82 = 'd0;
			end
			if (in_data164 < in_data165) begin
				temp_even83 = in_data164;
				in_data164 = in_data165;
				in_data165 = temp_even83;
			end
			else begin
				temp_even83 = 'd0;
			end
			if (in_data166 < in_data167) begin
				temp_even84 = in_data166;
				in_data166 = in_data167;
				in_data167 = temp_even84;
			end
			else begin
				temp_even84 = 'd0;
			end
			if (in_data168 < in_data169) begin
				temp_even85 = in_data168;
				in_data168 = in_data169;
				in_data169 = temp_even85;
			end
			else begin
				temp_even85 = 'd0;
			end
			if (in_data170 < in_data171) begin
				temp_even86 = in_data170;
				in_data170 = in_data171;
				in_data171 = temp_even86;
			end
			else begin
				temp_even86 = 'd0;
			end
			if (in_data172 < in_data173) begin
				temp_even87 = in_data172;
				in_data172 = in_data173;
				in_data173 = temp_even87;
			end
			else begin
				temp_even87 = 'd0;
			end
			if (in_data174 < in_data175) begin
				temp_even88 = in_data174;
				in_data174 = in_data175;
				in_data175 = temp_even88;
			end
			else begin
				temp_even88 = 'd0;
			end
			if (in_data176 < in_data177) begin
				temp_even89 = in_data176;
				in_data176 = in_data177;
				in_data177 = temp_even89;
			end
			else begin
				temp_even89 = 'd0;
			end
			if (in_data178 < in_data179) begin
				temp_even90 = in_data178;
				in_data178 = in_data179;
				in_data179 = temp_even90;
			end
			else begin
				temp_even90 = 'd0;
			end
			if (in_data180 < in_data181) begin
				temp_even91 = in_data180;
				in_data180 = in_data181;
				in_data181 = temp_even91;
			end
			else begin
				temp_even91 = 'd0;
			end
			if (in_data182 < in_data183) begin
				temp_even92 = in_data182;
				in_data182 = in_data183;
				in_data183 = temp_even92;
			end
			else begin
				temp_even92 = 'd0;
			end
			if (in_data184 < in_data185) begin
				temp_even93 = in_data184;
				in_data184 = in_data185;
				in_data185 = temp_even93;
			end
			else begin
				temp_even93 = 'd0;
			end
			if (in_data186 < in_data187) begin
				temp_even94 = in_data186;
				in_data186 = in_data187;
				in_data187 = temp_even94;
			end
			else begin
				temp_even94 = 'd0;
			end
			if (in_data188 < in_data189) begin
				temp_even95 = in_data188;
				in_data188 = in_data189;
				in_data189 = temp_even95;
			end
			else begin
				temp_even95 = 'd0;
			end
			if (in_data190 < in_data191) begin
				temp_even96 = in_data190;
				in_data190 = in_data191;
				in_data191 = temp_even96;
			end
			else begin
				temp_even96 = 'd0;
			end
			if (in_data192 < in_data193) begin
				temp_even97 = in_data192;
				in_data192 = in_data193;
				in_data193 = temp_even97;
			end
			else begin
				temp_even97 = 'd0;
			end
			if (in_data194 < in_data195) begin
				temp_even98 = in_data194;
				in_data194 = in_data195;
				in_data195 = temp_even98;
			end
			else begin
				temp_even98 = 'd0;
			end
			if (in_data196 < in_data197) begin
				temp_even99 = in_data196;
				in_data196 = in_data197;
				in_data197 = temp_even99;
			end
			else begin
				temp_even99 = 'd0;
			end
			if (in_data198 < in_data199) begin
				temp_even100 = in_data198;
				in_data198 = in_data199;
				in_data199 = temp_even100;
			end
			else begin
				temp_even100 = 'd0;
			end
			if (in_data200 < in_data201) begin
				temp_even101 = in_data200;
				in_data200 = in_data201;
				in_data201 = temp_even101;
			end
			else begin
				temp_even101 = 'd0;
			end
			if (in_data202 < in_data203) begin
				temp_even102 = in_data202;
				in_data202 = in_data203;
				in_data203 = temp_even102;
			end
			else begin
				temp_even102 = 'd0;
			end
			if (in_data204 < in_data205) begin
				temp_even103 = in_data204;
				in_data204 = in_data205;
				in_data205 = temp_even103;
			end
			else begin
				temp_even103 = 'd0;
			end
			if (in_data206 < in_data207) begin
				temp_even104 = in_data206;
				in_data206 = in_data207;
				in_data207 = temp_even104;
			end
			else begin
				temp_even104 = 'd0;
			end
			if (in_data208 < in_data209) begin
				temp_even105 = in_data208;
				in_data208 = in_data209;
				in_data209 = temp_even105;
			end
			else begin
				temp_even105 = 'd0;
			end
			if (in_data210 < in_data211) begin
				temp_even106 = in_data210;
				in_data210 = in_data211;
				in_data211 = temp_even106;
			end
			else begin
				temp_even106 = 'd0;
			end
			if (in_data212 < in_data213) begin
				temp_even107 = in_data212;
				in_data212 = in_data213;
				in_data213 = temp_even107;
			end
			else begin
				temp_even107 = 'd0;
			end
			if (in_data214 < in_data215) begin
				temp_even108 = in_data214;
				in_data214 = in_data215;
				in_data215 = temp_even108;
			end
			else begin
				temp_even108 = 'd0;
			end
			if (in_data216 < in_data217) begin
				temp_even109 = in_data216;
				in_data216 = in_data217;
				in_data217 = temp_even109;
			end
			else begin
				temp_even109 = 'd0;
			end
			if (in_data218 < in_data219) begin
				temp_even110 = in_data218;
				in_data218 = in_data219;
				in_data219 = temp_even110;
			end
			else begin
				temp_even110 = 'd0;
			end
			if (in_data220 < in_data221) begin
				temp_even111 = in_data220;
				in_data220 = in_data221;
				in_data221 = temp_even111;
			end
			else begin
				temp_even111 = 'd0;
			end
			if (in_data222 < in_data223) begin
				temp_even112 = in_data222;
				in_data222 = in_data223;
				in_data223 = temp_even112;
			end
			else begin
				temp_even112 = 'd0;
			end
			if (in_data224 < in_data225) begin
				temp_even113 = in_data224;
				in_data224 = in_data225;
				in_data225 = temp_even113;
			end
			else begin
				temp_even113 = 'd0;
			end
			if (in_data226 < in_data227) begin
				temp_even114 = in_data226;
				in_data226 = in_data227;
				in_data227 = temp_even114;
			end
			else begin
				temp_even114 = 'd0;
			end
			if (in_data228 < in_data229) begin
				temp_even115 = in_data228;
				in_data228 = in_data229;
				in_data229 = temp_even115;
			end
			else begin
				temp_even115 = 'd0;
			end
			if (in_data230 < in_data231) begin
				temp_even116 = in_data230;
				in_data230 = in_data231;
				in_data231 = temp_even116;
			end
			else begin
				temp_even116 = 'd0;
			end
			if (in_data232 < in_data233) begin
				temp_even117 = in_data232;
				in_data232 = in_data233;
				in_data233 = temp_even117;
			end
			else begin
				temp_even117 = 'd0;
			end
			if (in_data234 < in_data235) begin
				temp_even118 = in_data234;
				in_data234 = in_data235;
				in_data235 = temp_even118;
			end
			else begin
				temp_even118 = 'd0;
			end
			if (in_data236 < in_data237) begin
				temp_even119 = in_data236;
				in_data236 = in_data237;
				in_data237 = temp_even119;
			end
			else begin
				temp_even119 = 'd0;
			end
			if (in_data238 < in_data239) begin
				temp_even120 = in_data238;
				in_data238 = in_data239;
				in_data239 = temp_even120;
			end
			else begin
				temp_even120 = 'd0;
			end
			if (in_data240 < in_data241) begin
				temp_even121 = in_data240;
				in_data240 = in_data241;
				in_data241 = temp_even121;
			end
			else begin
				temp_even121 = 'd0;
			end
			if (in_data242 < in_data243) begin
				temp_even122 = in_data242;
				in_data242 = in_data243;
				in_data243 = temp_even122;
			end
			else begin
				temp_even122 = 'd0;
			end
			if (in_data244 < in_data245) begin
				temp_even123 = in_data244;
				in_data244 = in_data245;
				in_data245 = temp_even123;
			end
			else begin
				temp_even123 = 'd0;
			end
			if (in_data246 < in_data247) begin
				temp_even124 = in_data246;
				in_data246 = in_data247;
				in_data247 = temp_even124;
			end
			else begin
				temp_even124 = 'd0;
			end
			if (in_data248 < in_data249) begin
				temp_even125 = in_data248;
				in_data248 = in_data249;
				in_data249 = temp_even125;
			end
			else begin
				temp_even125 = 'd0;
			end
			if (in_data250 < in_data251) begin
				temp_even126 = in_data250;
				in_data250 = in_data251;
				in_data251 = temp_even126;
			end
			else begin
				temp_even126 = 'd0;
			end
			if (in_data252 < in_data253) begin
				temp_even127 = in_data252;
				in_data252 = in_data253;
				in_data253 = temp_even127;
			end
			else begin
				temp_even127 = 'd0;
			end
			if (in_data254 < in_data255) begin
				temp_even128 = in_data254;
				in_data254 = in_data255;
				in_data255 = temp_even128;
			end
			else begin
				temp_even128 = 'd0;
			end
		end
	end
	else begin
		temp_odd1   = 'd0;
		temp_odd2   = 'd0;
		temp_odd3   = 'd0;
		temp_odd4   = 'd0;
		temp_odd5   = 'd0;
		temp_odd6   = 'd0;
		temp_odd7   = 'd0;
		temp_odd8   = 'd0;
		temp_odd9   = 'd0;
		temp_odd10  = 'd0;
		temp_odd11  = 'd0;
		temp_odd12  = 'd0;
		temp_odd13  = 'd0;
		temp_odd14  = 'd0;
		temp_odd15  = 'd0;
		temp_odd16  = 'd0;
		temp_odd17  = 'd0;
		temp_odd18  = 'd0;
		temp_odd19  = 'd0;
		temp_odd20  = 'd0;
		temp_odd21  = 'd0;
		temp_odd22  = 'd0;
		temp_odd23  = 'd0;
		temp_odd24  = 'd0;
		temp_odd25  = 'd0;
		temp_odd26  = 'd0;
		temp_odd27  = 'd0;
		temp_odd28  = 'd0;
		temp_odd29  = 'd0;
		temp_odd30  = 'd0;
		temp_odd31  = 'd0;
		temp_odd32  = 'd0;
		temp_odd33  = 'd0;
		temp_odd34  = 'd0;
		temp_odd35  = 'd0;
		temp_odd36  = 'd0;
		temp_odd37  = 'd0;
		temp_odd38  = 'd0;
		temp_odd39  = 'd0;
		temp_odd40  = 'd0;
		temp_odd41  = 'd0;
		temp_odd42  = 'd0;
		temp_odd43  = 'd0;
		temp_odd44  = 'd0;
		temp_odd45  = 'd0;
		temp_odd46  = 'd0;
		temp_odd47  = 'd0;
		temp_odd48  = 'd0;
		temp_odd49  = 'd0;
		temp_odd50  = 'd0;
		temp_odd51  = 'd0;
		temp_odd52  = 'd0;
		temp_odd53  = 'd0;
		temp_odd54  = 'd0;
		temp_odd55  = 'd0;
		temp_odd56  = 'd0;
		temp_odd57  = 'd0;
		temp_odd58  = 'd0;
		temp_odd59  = 'd0;
		temp_odd60  = 'd0;
		temp_odd61  = 'd0;
		temp_odd62  = 'd0;
		temp_odd63  = 'd0;
		temp_odd64  = 'd0;
		temp_odd65  = 'd0;
		temp_odd66  = 'd0;
		temp_odd67  = 'd0;
		temp_odd68  = 'd0;
		temp_odd69  = 'd0;
		temp_odd70  = 'd0;
		temp_odd71  = 'd0;
		temp_odd72  = 'd0;
		temp_odd73  = 'd0;
		temp_odd74  = 'd0;
		temp_odd75  = 'd0;
		temp_odd76  = 'd0;
		temp_odd77  = 'd0;
		temp_odd78  = 'd0;
		temp_odd79  = 'd0;
		temp_odd80  = 'd0;
		temp_odd81  = 'd0;
		temp_odd82  = 'd0;
		temp_odd83  = 'd0;
		temp_odd84  = 'd0;
		temp_odd85  = 'd0;
		temp_odd86  = 'd0;
		temp_odd87  = 'd0;
		temp_odd88  = 'd0;
		temp_odd89  = 'd0;
		temp_odd90  = 'd0;
		temp_odd91  = 'd0;
		temp_odd92  = 'd0;
		temp_odd93  = 'd0;
		temp_odd94  = 'd0;
		temp_odd95  = 'd0;
		temp_odd96  = 'd0;
		temp_odd97  = 'd0;
		temp_odd98  = 'd0;
		temp_odd99  = 'd0;
		temp_odd100 = 'd0;
		temp_odd101 = 'd0;
		temp_odd102 = 'd0;
		temp_odd103 = 'd0;
		temp_odd104 = 'd0;
		temp_odd105 = 'd0;
		temp_odd106 = 'd0;
		temp_odd107 = 'd0;
		temp_odd108 = 'd0;
		temp_odd109 = 'd0;
		temp_odd110 = 'd0;
		temp_odd111 = 'd0;
		temp_odd112 = 'd0;
		temp_odd113 = 'd0;
		temp_odd114 = 'd0;
		temp_odd115 = 'd0;
		temp_odd116 = 'd0;
		temp_odd117 = 'd0;
		temp_odd118 = 'd0;
		temp_odd119 = 'd0;
		temp_odd120 = 'd0;
		temp_odd121 = 'd0;
		temp_odd122 = 'd0;
		temp_odd123 = 'd0;
		temp_odd124 = 'd0;
		temp_odd125 = 'd0;
		temp_odd126 = 'd0;
		temp_odd127 = 'd0;

		temp_even1	 = 'd0;
		temp_even2	 = 'd0;
		temp_even3	 = 'd0;
		temp_even4	 = 'd0;
		temp_even5	 = 'd0;
		temp_even6	 = 'd0;
		temp_even7	 = 'd0;
		temp_even8	 = 'd0;
		temp_even9	 = 'd0;
		temp_even10  = 'd0;
		temp_even11  = 'd0;
		temp_even12  = 'd0;
		temp_even13  = 'd0;
		temp_even14  = 'd0;
		temp_even15  = 'd0;
		temp_even16  = 'd0;
		temp_even17  = 'd0;
		temp_even18  = 'd0;
		temp_even19  = 'd0;
		temp_even20  = 'd0;
		temp_even21  = 'd0;
		temp_even22  = 'd0;
		temp_even23  = 'd0;
		temp_even24  = 'd0;
		temp_even25  = 'd0;
		temp_even26  = 'd0;
		temp_even27  = 'd0;
		temp_even28  = 'd0;
		temp_even29  = 'd0;
		temp_even30  = 'd0;
		temp_even31  = 'd0;
		temp_even32  = 'd0;
		temp_even33  = 'd0;
		temp_even34  = 'd0;
		temp_even35  = 'd0;
		temp_even36  = 'd0;
		temp_even37  = 'd0;
		temp_even38  = 'd0;
		temp_even39  = 'd0;
		temp_even40  = 'd0;
		temp_even41  = 'd0;
		temp_even42  = 'd0;
		temp_even43  = 'd0;
		temp_even44  = 'd0;
		temp_even45  = 'd0;
		temp_even46  = 'd0;
		temp_even47  = 'd0;
		temp_even48  = 'd0;
		temp_even49  = 'd0;
		temp_even50  = 'd0;
		temp_even51  = 'd0;
		temp_even52  = 'd0;
		temp_even53  = 'd0;
		temp_even54  = 'd0;
		temp_even55  = 'd0;
		temp_even56  = 'd0;
		temp_even57  = 'd0;
		temp_even58  = 'd0;
		temp_even59  = 'd0;
		temp_even60  = 'd0;
		temp_even61  = 'd0;
		temp_even62  = 'd0;
		temp_even63  = 'd0;
		temp_even64  = 'd0;
		temp_even65  = 'd0;
		temp_even66  = 'd0;
		temp_even67  = 'd0;
		temp_even68  = 'd0;
		temp_even69  = 'd0;
		temp_even70  = 'd0;
		temp_even71  = 'd0;
		temp_even72  = 'd0;
		temp_even73  = 'd0;
		temp_even74  = 'd0;
		temp_even75  = 'd0;
		temp_even76  = 'd0;
		temp_even77  = 'd0;
		temp_even78  = 'd0;
		temp_even79  = 'd0;
		temp_even80  = 'd0;
		temp_even81  = 'd0;
		temp_even82  = 'd0;
		temp_even83  = 'd0;
		temp_even84  = 'd0;
		temp_even85  = 'd0;
		temp_even86  = 'd0;
		temp_even87  = 'd0;
		temp_even88  = 'd0;
		temp_even89  = 'd0;
		temp_even90  = 'd0;
		temp_even91  = 'd0;
		temp_even92  = 'd0;
		temp_even93  = 'd0;
		temp_even94  = 'd0;
		temp_even95  = 'd0;
		temp_even96  = 'd0;
		temp_even97  = 'd0;
		temp_even98  = 'd0;
		temp_even99  = 'd0;
		temp_even100 = 'd0;
		temp_even101 = 'd0;
		temp_even102 = 'd0;
		temp_even103 = 'd0;
		temp_even104 = 'd0;
		temp_even105 = 'd0;
		temp_even106 = 'd0;
		temp_even107 = 'd0;
		temp_even108 = 'd0;
		temp_even109 = 'd0;
		temp_even110 = 'd0;
		temp_even111 = 'd0;
		temp_even112 = 'd0;
		temp_even113 = 'd0;
		temp_even114 = 'd0;
		temp_even115 = 'd0;
		temp_even116 = 'd0;
		temp_even117 = 'd0;
		temp_even118 = 'd0;
		temp_even119 = 'd0;
		temp_even120 = 'd0;
		temp_even121 = 'd0;
		temp_even122 = 'd0;
		temp_even123 = 'd0;
		temp_even124 = 'd0;
		temp_even125 = 'd0;
		temp_even126 = 'd0;
		temp_even127 = 'd0;
		temp_even128 = 'd0;
	end
end

endmodule